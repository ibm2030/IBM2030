-- CCROS library
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE std.textio.all;

package CCROS is
subtype CCROS_Address_Type is integer range 0 to 4095;
subtype CCROS_Word_Type is std_logic_vector(0 to 54);
type CCROS_Type is array(CCROS_Address_Type) of CCROS_Word_Type;
impure function readCCROS return CCROS_Type;
constant Package_CCROS : CCROS_Type :=
(
-- Replace below these comments, to the next comment
--          PCCCCCCPPCCCCCCCCCCCCCCCCCCCCCCCPPCCCCCCCCCCCCCCCCCCAAA
--          NNNNNNNSAHHHHLLLLMMMUUAAAABBKKKKKCDDDDFFFGGVVCCCSSSSASK
16#102# => "1111100110001000111001000000001011011000000000000000000",
16#10c# => "1000000000000111100000011100000000101011100000000000000",
16#169# => "1000011000000101100100011100001001011100100000000000001",
16#107# => "0011010111000000111001010011010000011001110010100000000",
16#181# => "0000001000001000100000011100000001111101100000000000000",
16#105# => "0100000100000000111001000000000111100100000000000000000",
16#1f3# => "0000001100000000100000011100000000111001100000000000000",
16#103# => "1111100000001000111001000000001011011000000000000000000",
16#1b6# => "1100010010001000011001000000000001000000000000000000000",
16#123# => "1101101011011000000100111100000001111101100001101010000",
16#109# => "0111000100010000000010011100001000101001100000000010000",
16#101# => "0000100010001000100100010000101000100001100000000000101",
16#1b4# => "1010001000001000100100000011011000100100001000000000000",
16#121# => "1101101101011000000100111100000001111101100001100000000",
16#116# => "0001000111000000100100111001000000111001111001010000000",
16#10b# => "1000101110001000000000000000000001101000000000000000000",
16#100# => "0000010001001000101100111011000101111001101000111100000",
16#2ec# => "1010001010001000100010000000000100100100000000011010000",
16#2e8# => "0111011001111111011001100000101110110011000000010000000",
16#2e4# => "1111010001110110100000100100010101100001111000110001001",
16#2e0# => "1111001011101110001100111000000000111001100001010110000",
16#2ed# => "0111000100000000100000100011001100101101001000000000000",
16#2e2# => "1111001100000000101100111000000001111001100001011011000",
16#2ee# => "1010001100001000100010000000000100100100000000011010000",
16#2ef# => "1110110010000100000000100000000000100101010000101001000",
16#200# => "1111010001110110100100111100000000111101100000010000000",
16#128# => "0000001000001000010001110011001101110001001000000000000",
16#2e9# => "1001010111111111000110100000000100110011000011010000000",
16#12a# => "1010100110001100000100110011001100110001001000000100000",
16#129# => "0111011010000000110001100000000001101101000000000000000",
16#12b# => "0111011100000000110001100000000001101101000000000000000",
16#131# => "0001011010001000000000111000000000111001100001010000000",
16#134# => "0001011010001101000100100111001100101111001000000111000",
16#133# => "0001101001100000000000111000000000111001100001010000000",
16#12c# => "1001100011010000101100011100000001110100100000000110000",
16#117# => "1000101100000000100100111100000000111101100000010000000",
16#2e5# => "1000101110110000100010100100000100100101111000110001000",
16#136# => "1011000100000100100100011100000001110001100000000000000",
16#137# => "0001101010001000000100110000000000111001100000000000000",
16#108# => "0001101011010000100000100000000000111101100001000000000",
16#12d# => "0000010000000000001100011100000001110100100000000110000",
16#184# => "0001011100000101100000011111001101101101001000000010000",
16#115# => "1100001111001000001100111000000000111001100000010111000",
16#2e7# => "1000101000110000100010100100000100100101111000110001000",
16#135# => "0001011100001000000100110000000000111001100000000000000",
16#186# => "1010001010001000100000000011010100100100001000001010000",
16#132# => "0001110010000000010101011100000001100001100001101011000",
16#140# => "1001100110001000000000100111001101101111001000000000000",
16#13d# => "0010000010000101010101110100000001110101111001100100000",
16#13c# => "1001111000111000100000101100000001101101100010000110000",
16#10a# => "1001111101011000010101110000000000110001111001000000000",
16#138# => "0000010010001000000000101100000001101101100010000000000",
16#12e# => "0001110100000100110101011100000001110001100000000000000",
16#141# => "1010010001101110100000011100000000100001100001101001000",
16#13f# => "0010000000000000110101110100000001110101111001100100000",
16#139# => "0001110000000000000100111100000000111101100000010000000",
16#145# => "1010010111101110100000100000000000100001111001101001000",
16#144# => "1010001000000000110101110100000001110101111001100100000",
16#13e# => "1010001111100000000000101100000001101101100010000000000",
16#13a# => "1010010001101110100100000000000000100000000000000110000",
16#12f# => "0001110110001100100100011100000000110001100000000100000",
16#13b# => "0001110010001000000100111100000000111101100000010000000",
16#30d# => "1010001000001000100110000000000100100100000000011010000",
16#385# => "1000011100010000100000100010000000101100101000000000000",
16#375# => "1100001000000000111001100101110001100000101000000010000",
16#30f# => "0111101110001001000100001101000001101000010000010000100",
16#39c# => "1111100010000100010001100011001100101101001000000000000",
16#2eb# => "1100111001111111000110100011001110110011001001000100000",
16#388# => "1000000011000111101010000000000100100100000000001000000",
16#3cc# => "1100010110000000011001100100110000011101100000001010000",
16#39e# => "1111100000001100010001100011001100101101001000000000000",
16#39f# => "1111100110001100010001100011001101101101001000001011000",
16#397# => "0000001100000000000110101111000100000011111000100001000",
16#39d# => "0100101100001000100100100011001100101101001000000000000",
16#2d4# => "1001001000000000000110000000000101000000000000000000000",
16#2da# => "1110101110000000000000100011001100101101001000000000000",
16#2ea# => "1110110010001111011001100000110000110011000000010000000",
16#125# => "1010001110001000100100000000000000100100000000011010000",
16#2db# => "1001001100010000100010101011000100101001110000110000000",
16#127# => "0111101101000000111001111000001011011101100000001011000",
16#142# => "1000000101000111101000000000000000100100000000001000000",
16#190# => "0010000100001000010000000000000001000000000000001010000",
16#15d# => "1100100111001101100000110000000001110001100001100000000",
16#154# => "1010111011011000110101101100000001101101100011001101000",
16#182# => "0010101001111100000000100111001100101101001000000110000",
16#14c# => "0100000010001111011001100000000001011101100000001011000",
16#148# => "0010011101110011100100110011000101000001101000101001000",
16#192# => "0010000010001000010000000000000001000000000000001010000",
16#15f# => "1010001100001000100000000011010100100100001000001010000",
16#156# => "1010111001011000110101000000000000000000000001001100000",
16#14d# => "0100000000001111000100000000000001000000000000001010000",
16#143# => "0010101010001000001000000000000001000000000000000000000",
16#191# => "0010000110001000110000110000000000110001100010000000000",
16#15e# => "1010001010001000100000000011010100100100001000001010000",
16#157# => "1010111011011000010000000000000001000000000000000000000",
16#185# => "0010000010001000010101000000000001000000000000001010000",
16#15c# => "1100001000000000100000000000000001000000000000000000000",
16#183# => "0010110011111100001000100111001101101101001001000110000",
16#197# => "0010000010001000010101000000000000011100000000000110000",
16#193# => "1010001000001000100100000011011000100100001000001010000",
16#14e# => "1010001000001000100100000011010100100100001000001010000",
16#194# => "0100101110001000010101110100000001011101100000001101000",
16#196# => "0100101100111101101000101100000001101101100010001010000",
16#155# => "0100101100001000010101110000000000011101100000001100000",
16#3c2# => "1010001100001001000100000111011000100100001000001010000",
16#14f# => "1110000011001111000110100111001110101101001000001010000",
16#195# => "0100101000001000010101100000000001011101100000000111000",
16#3c3# => "1010001010001001000100000111011000100100001000001010000",
16#1a3# => "1010001100001000100000000000000000100100000000011010000",
16#18c# => "1010001110001000100100000011010100100100001000001010000",
16#149# => "0100011010011011100100110011001101110001101000001011000",
16#1a2# => "1010001010001000100000000000000000100100000000011010000",
16#18d# => "1010001000001000100100000011011000100100001000001010000",
16#1a1# => "1010001010001000100000000000000000100100000000011010000",
16#18e# => "1010001000001000100100000011010100100100001000001010000",
16#1a0# => "0000111000000000010101000000000000100100000000001101000",
16#198# => "1101000111111100000000000000000000000000000000000100000",
16#18f# => "0100110111110111010011100111001100101101001000001100000",
16#19b# => "1100111011111000000000101111000100000011111000100001000",
16#318# => "1001001011111111000100100111001100101101001000001010000",
16#164# => "1000110111110110100010011100001110100001100001101001000",
16#146# => "0011001111101110010101110100000000110101111001100000000",
16#166# => "1010001100001000100000000000000000100100000000011010000",
16#3f6# => "1010001010001001000100000111010100100100001000001010000",
16#319# => "0111101101001111000100100100000001101101000000000000000",
16#160# => "0011001101101110000100000000000001011100000001000000000",
16#3f7# => "1010001100001001000100000111010100100100001000001010000",
16#161# => "1011000110000000000100111100000000111101100000010000000",
16#31e# => "1010001010001001000100000111010100100100001000001010000",
16#31b# => "0000111111001111000100101011010000101110110000011001000",
16#165# => "0011100001000101100010011100001110101101100001101001000",
16#167# => "0011100111000101100010011100001111000001100001101001000",
16#371# => "0000001110001000000000111100000000111101100010000000000",
16#3a1# => "0011100000000000100100111100110000011101100000000000001",
16#376# => "1000101100000000101010111100000100111101100000001101000",
16#32a# => "1011101000001000011001101011010001011110110000000000000",
16#306# => "1001010110001000000000010011010000011001110000110000000",
16#3a0# => "0000001110001000000100111100110000011101100000000000001",
16#35f# => "1101000110000100111001111100000111111101100001100000000",
16#384# => "1010111110001000101000110100001100100001100000000000001",
16#370# => "1100001100000000011001111011001010011101101001000000000",
16#374# => "1010001010001001000100000111010100100100001000001010000",
16#35d# => "1011101100000000000100000011010000101000010000000000000",
16#3f8# => "1010001100001001000100000100000000100100000000011010000",
16#372# => "1011101010001000000100110100001100100001100000000000001",
16#37d# => "1010001010001001000100000100000000100100000000011010000",
16#30e# => "1000011000000000000100111100000000111101100000010000000",
16#38b# => "1010001010001001000100000111010100100100001000001010000",
16#3fa# => "1010001010001001000100000100000000100100000000011010000",
16#30c# => "0011111011110111000100110100000000110101100001100000000",
16#389# => "1000011100110000000100110001000001110001101001000000000",
16#3fb# => "1100010101001000100100111010000001111001101000000000000",
16#373# => "0111110001101110100100100100000000100011100000000010000",
16#3f9# => "1000101011110111000100101100000001000001100000000110000",
16#168# => "1000000110000000001000110000000000111001100000000000000",
16#1a8# => "0011010010000000011001101011010001011110110000000000000",
16#1a7# => "0101010110000000001000010011010000011001110000110000000",
16#1a5# => "0101001100001000111001111000001010011101100000000000000",
16#1a4# => "0101001010000000101000110100110001111101100000000000001",
16#19d# => "0101001111010000011001111100000110011101100000000000000",
16#187# => "1100111001000000100000011100000001100101100000000000000",
16#158# => "1100001010001000110101101100000001000001000000000010000",
16#1a6# => "0101001000000000001000000000000001100100000000000000000",
16#19f# => "1010001000001000100100000011001100100100001000001010000",
16#272# => "0011100100000101000000110000000001110001100000011000000",
16#2d8# => "0011100100001000010001100011001100101101001000000000000",
16#214# => "1000000001000111100010000000000101011000000000000000000",
16#2d9# => "1000101111001101010001110011001001110001101000001000000",
16#281# => "1000000000000111100010011100000101111101100000000110000",
16#201# => "0100000011000000110001111011000101100101101000101001000",
16#284# => "1000000100000000101000000000000001000000000000000000000",
16#203# => "1100001000000000011001100100000001011101100000001011000",
16#215# => "1000000111000111100010000000000101011000000000000000000",
16#283# => "0000111110001000100000011100000000110101100000000000000",
16#2c1# => "1000000011001000100000011100000000111001100000000000000",
16#206# => "1110000000000000110001110000000000110001100010000000000",
16#216# => "0000001010001000000000011100000001100101100000001001000",
16#275# => "1000000011000111100110000000000101011000000000000000000",
16#217# => "1000000001000111100010000000000100100100000000001000000",
16#221# => "0000111000000000100100000011010000101000010000000000000",
16#261# => "0001000010000000101000010011010000011001110010100000000",
16#21f# => "1011000110000000111001000000010000011100000000000000000",
16#277# => "1000000101000111100110000000000101011000000000000000000",
16#2fd# => "1011101011001011100100000000000001100100000000000000000",
16#1aa# => "1111111000000000100010011101001000000001010000100000000",
16#15b# => "0101010010001000011001000000101111000000000000000000000",
16#21d# => "1000000100000111100110110100000101111101100000000110000",
16#274# => "0000111001000000100100110000000000111001100000000000000",
16#276# => "1011101010000000000100110011000101100101101000100000000",
16#271# => "0000001100001000110101110011000101000001101000101001000",
16#280# => "0011100010000000101000000000000000000000000000001011000",
16#273# => "0100000110000000011001100100000000011101100000000000000",
16#205# => "0011100101001000100000011100000001110001100000000000000",
16#204# => "0000001010000000110001011100000000110101100000000000000",
16#202# => "0000001010000000000000110000000000110001100000010000000",
16#270# => "1000000010001000010001011100000001100101100000001001000",
16#211# => "1011101101001101000000000000000001100100000000000000000",
16#20c# => "0000100100000100110101101100000001000000100000000111000",
16#208# => "1000011010000011100000101100000001101101100010000000000",
16#207# => "0000010010000000000100011100000000011101100011000000000",
16#15a# => "0000001100001001010101001000000001000000000000000110000",
16#20b# => "1011101011001101000000000000000001100100000000000000000",
16#210# => "0000010010111011100100011100000001011101100011100000000",
16#20d# => "0000100010000000010101101100000000000000100000000000000",
16#20a# => "1000011100000011100000101100000001101101100010000000000",
16#20e# => "1011101111001101000100000000000001000000000000000000000",
16#209# => "1000011100001011100000000000000001100100000000000000000",
16#20f# => "1000000101000111100110000000000101011000000000000000000",
16#2dc# => "1010100010000000100010101100000011101101000000000000000",
16#1b1# => "1101011101000000101000110011000101000001101000101001000",
16#1b2# => "0101100101001000100000011100000001110001100000000000000",
16#1b0# => "0101100010001000010001011100000001110101100000000100000",
16#130# => "0101100100000000000000110000000000110001100000011010000",
16#1ac# => "1001100000000000010001011100000001100101100000001001000",
16#2dd# => "1101011001000101000010110000000101110001100000011000000",
16#2e1# => "0110111100000100010001011100000001100011100000000000000",
16#1b3# => "0101100010000000111001100100000001011101100000001011000",
16#1ae# => "1001100110000000010001011100000001100101100000001001000",
16#1ad# => "0011010110001000010101111000000000011101100000000000000",
16#1af# => "1111100000001000111001000000001011000000000000000000000",
16#33d# => "1011101001001000000010011100001001110001100000000000000",
16#33a# => "1001111110110100011001000000101011100100000000000000000",
16#337# => "0001110000001011000100101001000000100101110001100000000",
16#329# => "0001011100001000000100100111001100110011001000001100000",
16#32c# => "1001010001001000101000110011000101000001101000101001000",
16#327# => "0001011010000000011001110000101010011101100011010100000",
16#33e# => "1011101001001000000010011100001001110001100000000000000",
16#386# => "0001011100001000001000100111001100110011001000001100000",
16#32b# => "1100001110001000011001100000000001011101100000001011000",
16#33c# => "1000000111000111100010000000000101011000000000000000000",
16#33b# => "1001111001100100011001000000101011100100000000000000000",
16#33f# => "1000000111000111100010000000000101011000000000000000000",
16#32e# => "1001100110000000010001110011000100000001110000100010000",
16#339# => "0001101010001000100000100100000000100101111011100000000",
16#334# => "0001110000000101000100011110000000011101111000000000000",
16#336# => "0001101110000101110101011100000001100101100000000000000",
16#331# => "0001101000001000000000110000000000110001100010000000000",
16#332# => "1001100101010000110001011100000000100001100000000000000",
16#330# => "1001100010001000000000110011000100110001110000110000000",
16#32d# => "1001100010000000010001100100000000100101111011101100000",
16#338# => "0001011100110000100000101100000000101101100010000001000",
16#335# => "0001110110000101000100011110000001011101111000010000000",
16#333# => "0001101010001000000000110011000101110001111010010000000",
16#32f# => "1001100100000000010001100100000001100101111011101101000",
16#124# => "1101110001111100011001100000100100100101100000000100000",
16#1bb# => "1010001100001000100000000000000000100100000000011010000",
16#1c2# => "1010001010001000100000000011011000100100001000001010000",
16#1be# => "1010001100001000100000000011010100100100001000001010000",
16#1bc# => "1010001110001000100000000011001000100100001000001010000",
16#1b8# => "1101101000000000100000011111111001100101101010100001000",
16#1c3# => "0110001100000100000000011100000001110101100000000111000",
16#1c0# => "1110000000001011110001011100000001110001100000000000000",
16#1bf# => "1110000110000000000000011100000000000000100000000000000",
16#1b7# => "0101111100001011110001110000000000110001100010000000000",
16#1bd# => "1101101000001000100000011100000001000001100000000000000",
16#1b5# => "0101111110000101010001110011001000110001101000000000000",
16#1b9# => "1101101110000000100000011111111001100101101010100001000",
16#1cb# => "0110001010000000100000011100000000100010100000000110000",
16#1c4# => "0110010010111000110101100000000000011101100000000000000",
16#1ca# => "0110001000000000000000010100000000100011000000000110100",
16#1c9# => "1000000101000111101000000000000000100100000000001000000",
16#1c8# => "0110010110000000100100100110000001001101001000000000000",
16#1c5# => "0110010100111000010000000000000001000000000000001010000",
16#3df# => "1010001100001000100010000000000100100100000000010000000",
16#48c# => "1001111011010010101000101100000000100001100000000000000",
16#48a# => "0100011011001000010101101100000000101101100000010010000",
16#489# => "1100010010001000000000011100000001000001100000001001000",
16#43d# => "1100010010000000110000110000000000110001100000010000000",
16#3d3# => "1001111000000000100110101100010000100001100000000000000",
16#48e# => "1001111001010010101000000000000001000000000000000000000",
16#492# => "0110001010000010100100100000000000110001100001000110000",
16#490# => "1100100100001011100100011100000001011101000000001010000",
16#48b# => "1100100100000011100100011111101101000000101010010000000",
16#43e# => "1100010110001000100100011111110100000000101010010100000",
16#494# => "0100110010000000000100100000000000110101100000000000000",
16#4c5# => "0100101000000000000100100111001100101101001000001100000",
16#493# => "0110001100000010100100100000000001110001100011010111000",
16#491# => "1100100010001000100100011100000001011101000000001010000",
16#43f# => "1010001000001001000100000111011100100100001000001010000",
16#43c# => "1010001000001001000100000111011100100100001000001010000",
16#4c4# => "1010001110001001000100000111011100100100001000001010000",
16#49c# => "1010001100001001000100000111100100100100001000001010000",
16#49f# => "1100111000000100100100000011100100100100001000001010000",
16#4da# => "1010001010001001000100000111100100100100001000001010000",
16#49d# => "1110110111001000000100000000000001100100000000000000000",
16#4d8# => "1000000101000111100110000000000101011000000000000000000",
16#49e# => "1110110111001000000100000000000001100100000000000000000",
16#449# => "1100111110111011100100110110000001000001110000011001000",
16#44a# => "0100101110000000110001100010000001100100101000000000000",
16#443# => "1010010111001000001000110000000000110001100000010000000",
16#442# => "0010000000001000110001100000000001011110110000001001000",
16#440# => "0010000010001000000100011110000000100000111000001101000",
16#448# => "1010010000001000000100110100000001110101100000010000000",
16#497# => "0010000010000101100100100001000000100001111000000000000",
16#496# => "0100101000001000100100100010000000100001111000000000000",
16#495# => "0100101000001011100000100101000000100001111000000000000",
16#4c7# => "0100101010000000100100100010000001100100101000000000000",
16#499# => "0110001100001010100100011110000000011100110000000000000",
16#441# => "0100110000000000100000011110000000100010111000001100000",
16#498# => "0010000110000000110001000000000001100000000000001000000",
16#4c2# => "0100110010001000101000101100000000101101100010000001000",
16#49a# => "1110000000001101010101000001000001011100011101100000000",
16#447# => "0100110000001000001000101001000001100100110000001010000",
16#4c6# => "1010001001011000110001100000000001100111000000000000000",
16#4c3# => "1010010100000000101000011111100000000001110000101000000",
16#49b# => "0100110010000000000100110100000001110001100000000000000",
16#445# => "0100110010001000101000101010000000101001001000001011000",
16#4a2# => "0101001010011101101000100100000001101101000000000000000",
16#4a4# => "1101000010001000010000110000000000110001100000010000000",
16#3d2# => "0101001110000000000110000000010000011100000000000000000",
16#4a5# => "1101000100001000010000110000000000110001100000010000000",
16#4a6# => "1101000100001000010000110000000001110001100000011101000",
16#4b7# => "0101010000000000100100101100000001101101100000010000000",
16#4b8# => "1101101001001000100000000000000001100000011010001001000",
16#4b0# => "1101110011010101010101101111001100000000101010010001000",
16#4a3# => "0101100100000000000000011111100001000001010000100010000",
16#4a7# => "1101000110001000110101110000000001100101100010000100000",
16#4b5# => "0101100011001000000100101100000001101101100000010000000",
16#4ba# => "1101101011001000100000011100000000100001100000001001000",
16#4b9# => "0000010010001000000000000000100101100000000011010110001",
16#4bb# => "0000010100001000000000000000100100100000000011000110001",
16#4b3# => "0101100010000000000100110011011100110001101000110000000",
16#4b4# => "1101011000001101101000100010000001100001111001101101000",
16#4ae# => "1101101010000000000100011100000000011101111111101010000",
16#4aa# => "1101011000001000000000100010000000100001111001101100000",
16#4a9# => "0101010100001000010000000000000000000000000010001001000",
16#4b2# => "0101010100000000100100110000000000110001100010000000000",
16#4b6# => "0101010011001000001000110001000000000000101010011000000",
16#4af# => "1101101001011000010000011100000001011101111111101011000",
16#4ac# => "0101010100000000100100110000000000110001100010000000000",
16#4a8# => "1101011010000011100100100010000000100001111001100000000",
16#4ad# => "0101100110001011100100100100000000100101100010001001000",
16#4bf# => "1000000011000111101010000000000101100100000000001010000",
16#4c0# => "0101111100001101010000101110000001011111001000000000000",
16#4bd# => "1110000000000000000000011100000001101101100111101000000",
16#4db# => "0101111000000000110000110001000000000000101010010001000",
16#408# => "1110110011001000100100100011101100100000101000000000000",
16#4be# => "1110110000000000101000101100000000100010100000000000000",
16#4d9# => "1110110110001000100100110000000000110001100010000000000",
16#40a# => "1110110101001000100100100011110100100000101000000000000",
16#704# => "1010001010001001000100000111011000100100001000001010000",
16#703# => "0000001100000011100000000011011100101100001010001010000",
16#700# => "1000000000001111010001110011000101000001110000100000000",
16#3ac# => "1000000110000000000110100100011101110001000011010000000",
16#31a# => "1101011000000000000100110011110001100001110010100000000",
16#705# => "0000001000001100000100011111100000000010101000100001000",
16#702# => "0000001110000000100000000011001101101100001010001011000",
16#70c# => "0010011101010100000110110000010001110001100001100110000",
16#70d# => "0010011011010100000110110000010001110001100001100110000",
16#70b# => "1000011111111101000100100010000000100101111000000010000",
16#708# => "0000010010001100000100101001000001101001110000001000000",
16#701# => "0000010010000000000100110111001101100111010000100000000",
16#707# => "1000000110000000100100100000000000110101100000000000000",
16#70e# => "0010011011010100000110110000010000110001100001100111000",
16#706# => "1000000000000000100100000010000000110100011010010000000",
16#70f# => "0010011101010100000110110000010001110001100001100110000",
16#70a# => "1000011001111101000100100010000000100101111001000011000",
16#460# => "0010011001010000100000110000000001110001100000011000000",
16#4e0# => "1011000111001000010001100111000101100101110010010010000",
16#44d# => "0111000100011111000100000000000000000000011100001001000",
16#462# => "1011000110000000000100000000000000000000000011010000000",
16#4e1# => "1011000001001000010001100111000101100101110010010010000",
16#4e3# => "0111000110000000100100110011000100110001010000001011000",
16#4ee# => "0111011000001000101000000000000000100100000011010000000",
16#4ef# => "0101100110001000000110101100001001101101100000011001000",
16#4ec# => "0111011010001101001000000000000001100100000000000000000",
16#4e2# => "0111011001001000010101000000000000011100000000000000000",
16#714# => "0011111101001000100110000000001000100100011100000000000",
16#710# => "1000101010011101100100011111011100000001101010101001000",
16#27f# => "0011111010000000100100000000000000000000000011010000000",
16#71e# => "0000100001101110100100000000000000100100000000001000000",
16#461# => "0000111110001011100110000000011101011100011100001100000",
16#44f# => "1011000010000000100100100011010001000001101000100000000",
16#715# => "0011111011001000100110110000001000110001100010000000000",
16#711# => "1000101000011101100100011111001100000001101010101001000",
16#71f# => "0000111110001000000100011100000001011110100000001101000",
16#717# => "0011111101001000100110110000001000110001100010000000000",
16#712# => "1000101100011101100100011111000100000001101010101001000",
16#293# => "1100100100000000100100000000000000000000000011010000000",
16#26c# => "0011111001001000100100110011000100110001010000001011000",
16#26e# => "1100100011001000100100100100000001011111000000001101000",
16#716# => "1011011011011000000110000000001000100100011100000000000",
16#713# => "1000101110011101100100011100000001000001100000001001000",
16#40d# => "0010011011010000001000101100000001101101100000010000000",
16#47d# => "1000011000000000110101100111000101100101110010010010000",
16#44c# => "0011111010110000100100000000000001011100000100000000000",
16#419# => "1111001110000000000100101011001101101001110010100100000",
16#47f# => "1000110010000000100100000000000001101100000010001010000",
16#2f8# => "1011000110001000010001110000000000110001100000011100000",
16#47e# => "1000110100000000100100000000000001101100000010001010000",
16#44e# => "0011111000110000000100100111100100000011010010010000000",
16#2f9# => "1011000000001000010001110000000001110001100000011101000",
16#47c# => "0111110110110101000110000000001000100100000100000000000",
16#2fa# => "1111100100000000100100000000000000011100000100001101000",
16#26d# => "1011011010001000100100110011000101110001010000000000000",
16#2f4# => "0111101010000000100100100100000000011111000000000000000",
16#269# => "0011001000000000101000101100000001101101100000010000000",
16#2f0# => "0011010100000000110101011101000001011110110000000000000",
16#262# => "1111100110011101100000100100000001100111001000001000000",
16#265# => "1011000100001011110001110000000000110001100000010000000",
16#26f# => "1111001001101100100110011100010001100101111001000100000",
16#2f5# => "1011011001011000100100000000000001101100000010000000000",
16#2f1# => "0011010010000000110101000000000001000000000000000000000",
16#27d# => "1011000000001000010001110000000000110001100000010000000",
16#2f6# => "0011111100001000010101100100000001011111000000001101000",
16#27c# => "0011010110000000101000110011000100110001010000001011000",
16#2f2# => "0011111011011000010101011101000001011110110000000000000",
16#2f7# => "0011111010001000010101000000000001000000000000000000000",
16#282# => "0111101101001101100100000000000001011100000000001000000",
16#27e# => "0100000000001000001000101100000001101101100000011001000",
16#2f3# => "0011111101011000010101000000000001000000000000000000000",
16#291# => "0011111010001000010101000000000000000000000000001000000",
16#263# => "0111101000000101100000000000000001000000000000000000000",
16#4e4# => "0011100100000000100100110011001100110001001000001000000",
16#478# => "0011100100110000100100110011001101110001001000001010000",
16#4a0# => "0011100100110000100100110011001101110001001000000000000",
16#4e5# => "1111001110000000000100000000000000000000000000000001000",
16#47a# => "0011100010110000100100110011001100110001001000001011000",
16#4a1# => "1011110010110000000100100101000001000001111000000000000",
16#4e6# => "1101000110000110100100100101000000100101111000001000000",
16#4e7# => "1111001100001000000100000000000000000000000000000001000",
16#4e8# => "1000000101000111100110000000000100100100000000001000000",
16#47b# => "0101010000001000100100011111100001011101110000111100000",
16#4e9# => "1000000011000111100110000000000100100100000000001000000",
16#4ab# => "1110110110000000100010000000000101000000000000000000000",
16#479# => "0101010110001000100100011111100001011101110010101100000",
16#4eb# => "1011110100111000110001000000000001000000000000000000000",
16#4ea# => "1110110110000000000110101000000100000001010000100000000",
16#48d# => "0011100100110000101000110000000000110001100010001010000",
16#470# => "0100011110000000110001100100000000011101100000001001000",
16#4f8# => "0011100110011000000000011100000001100101100000000000000",
16#471# => "0111110101101110110101101100000001101101100010001100000",
16#48f# => "0011100010110000101000110000000001110001100010001011000",
16#472# => "0111101000000111010001100100000000011101100000001001000",
16#4f9# => "0011100000011000000000011100000001100101111001100000000",
16#473# => "0111110011101110110101101100000000101101100010001101000",
16#4f0# => "0100011100110000110001100101000000011101111000001001000",
16#4fa# => "1111100100011101100000011100000001100101111001100000000",
16#409# => "0011100000000000100100101011010000101001101010101100000",
16#4f5# => "0000010100110000101000110011110001110001101010001010000",
16#4f1# => "0100011010110000110001100101000001011101111000011001000",
16#464# => "1111100110011101100100100101000001100101111000000000000",
16#4fb# => "0011001011011000000000011100000001100101111001100000000",
16#40b# => "0011100010001000100100101011010001101001101010101101000",
16#4f7# => "0000010010110000101000110011110000110001101010001011000",
16#4f2# => "0111101010110111010001100101000000011101111000001001000",
16#466# => "1111100000011101100100100101000000100101111000010000000",
16#4f4# => "1111010011111101001000000011100000101000010000001010000",
16#4f3# => "0111101100110111010001100101000001011101111000011001000",
16#4f6# => "1111010101111101001000000011100000101000010000001010000",
16#1d0# => "1110011110001000000000000000000001000000000000000000000",
16#3f0# => "0110001010001000100010000000000101100100000001001011000",
16#1c1# => "1101000110001110100010011100001110100001100000000000000",
16#1ce# => "1110000110000000110011101100000000101101100010000001000",
16#1d2# => "1110011000001000000000000000000001000000000000000000000",
16#3a4# => "0110100101011101000110011110000101011101111101101001000",
16#3a3# => "0101001010000101110101110000000000110001100010000000000",
16#3f1# => "1101000000001000100000011100000000100001100011011101000",
16#19a# => "1111100101111100000110000000001111000000000000001010000",
16#1cf# => "1110110000110011000100100011100000100001110000100000000",
16#3a5# => "1110011110001101000010011110000101100001111011101001000",
16#3a2# => "0101001000001101110101011111100000000001110000100010000",
16#3f2# => "1101000000001000100000011100000001100001100001000000000",
16#1d1# => "1110110100110011000000011111100001000001110000100000000",
16#1fc# => "1101011101010000100010101100001110101101100010000001000",
16#3a7# => "1111111000000101000110011110000101100001111011101001000",
16#3af# => "0101001110001101110101000000000000100000000000000000000",
16#3f3# => "1101000110001000100000011100000000100001100011010111000",
16#19e# => "1111100110001100000110000000001110000000000000000100000",
16#1fd# => "1110110010110011000000100011100000100001110000100000000",
16#3ab# => "1111100101111100010011000000000001000000000000001010000",
16#3c0# => "0101010110001000100100110000000000110001100000011100000",
16#1d5# => "1110110010110011000000011111100000100001110000100000000",
16#1d3# => "0111000011001100100000000000000001000000000000000110000",
16#1d4# => "1101011101010000100010101100001110101101100010000001000",
16#3a6# => "1110101110000101000110011110000101011101111101101001000",
16#3ad# => "0101001000001101110101010011111100100001111000000000100",
16#1e8# => "1111001100000000100100011111100000011100110000001010000",
16#1e9# => "1111001010000000100100011111100000011100110000001010000",
16#1e0# => "1111010010000000111001000000101111000000000000000000000",
16#1ea# => "1111001010000000100100011111010000011100110000001010000",
16#1e2# => "1111010100001000011001000000101111000000000000000000000",
16#1d8# => "1111010101001011111001000000101111000000000000000110000",
16#1eb# => "1111001100000000100100011111001000011100110000001010000",
16#1e1# => "1111010000001000111001000000101111000000000000000000000",
16#1db# => "1111010101001011111001000000101111000000000000000110000",
16#1e5# => "1000000011000111101000000000000000100100000000001000000",
16#1df# => "1111001010000000100100011111000100011100110000001010000",
16#1e3# => "0110111110001000111001000000101111000000000000000000000",
16#1d7# => "1110110100001000100000100011100001000001110001110000000",
16#1d9# => "1110101110001101111001000000101110100100000000010000000",
16#1e4# => "1010001100001000101000000011100001100100001000001000000",
16#1dd# => "1111001100000011111001100100101111011111001000001010000",
16#1d6# => "0110111110000000100000011111100000000000101000100110000",
16#1da# => "1110101110001101111001000000101110100100000000010000000",
16#1ec# => "0011100010001000000000011100000001100101100000000000000",
16#170# => "0111011110000011110011101100000001101101100000010000000",
16#396# => "0011100010011000000010000000000100000000000001000000000",
16#398# => "0100101100001000000100011101000001011101111000101001000",
16#387# => "0100110011111100010101110000000000110001100000010000000",
16#1ed# => "1100001000001000100010011100001111100101100000000000000",
16#1e6# => "0111011110000000110011101100000001101101000000000000000",
16#199# => "1111001000001000000000110011001100110001101010100000000",
16#39a# => "0100101010001000000100011101000000011101111000111001000",
16#3f5# => "0100110011111100010000000000000001110000000000000000000",
16#39b# => "0100101100001000000100011101000001011101111001111001000",
16#172# => "1111010001001100111001000000101111000000000000000110000",
16#399# => "0011100010011000000010011101000100000001111011011001000",
16#119# => "1011101010001000010101000000000001000000000000000000000",
16#11a# => "1011101010001000010101000000000001000000000000000000000",
16#11b# => "1011101100001000010101000000000000011100011011010111000",
16#118# => "1011101100001000010101000000000000011100011011010111000",
16#1ee# => "1000110101010100000000011100000001000001100000001001000",
16#10e# => "0111011110001000010001011111100000000001110000100010000",
16#106# => "1000011100001000000000100011001101101101001001000000000",
16#176# => "1010100010000101101000110000000000110001100010000000000",
16#1ef# => "1011101110001101010000101100000000101101100010000001000",
16#11c# => "0111011010001000100000000000000001000000000000000000000",
16#151# => "0000111110000000010101000000000001000000000000000000000",
16#174# => "1010100000000000001000110000000000110001100010000000000",
16#1c7# => "1011101011011101010101000000000001011100011101101001000",
16#11d# => "0110001100001110100000000000000001000000000000000000000",
16#150# => "0000111000000000110011101100000000101101100010000001000",
16#175# => "1110110110110011001000011111100001000001110000100000000",
16#1c6# => "1110011000000000010101011111100000000001110000100010000",
16#152# => "0000111010000000110001100011001101101101001001000000000",
16#177# => "1000000101000111101000000000000001011000000000000000000",
16#1cc# => "0110111101010000001000101100000000101101100010000001000",
16#1de# => "1110011000000101010101000000000000011100000000000000000",
16#153# => "0000111100000000110001100011001101101101001000000111000",
16#1cd# => "1000000011000111101000000000000001011000000000000000000",
16#1dc# => "1110011110000101010101000000000001011100000010000000000",
16#38c# => "1010001100011000000000000000000000000000000010001001000",
16#38e# => "1000000011000111101010000000000101100100000000001010000",
16#3f4# => "0100011101111100010000100100000001011101100000001101000",
16#392# => "0100011000001000011001100000101110011101100000000000000",
16#390# => "1100100010001011100000011111010000100000110000000000000",
16#345# => "1100100100000011111001100001101110000001111001110000000",
16#38d# => "1010001110000000100000100100000001100001111000100000000",
16#393# => "0100011010001000011001101000101111011111001000000000000",
16#391# => "0100011100001000000100011111100000011100110000000000000",
16#3c5# => "0011100110001000000010000000000100000000000000001000000",
16#38f# => "0110001000010000100100000000000000011100000011001001000",
16#3c7# => "0011100000001000000010000000000101000000000000000000000",
16#347# => "1010001110001000000100110100000001110101100000010000000",
16#394# => "1010001100001100100000101111001100000000101001111001000",
16#34c# => "0100101100000101110000110000000001110001100001010000000",
16#34a# => "0010011100000000001000101100000001101101100000010000000",
16#346# => "1010010101001101110101101101000000000010101001111000000",
16#3fc# => "1010001010011000000000110000000001110001100001011100000",
16#31c# => "1111111101111100010000100100000001101101000000000000000",
16#395# => "1010001110001100101000101111001100000000101001111001000",
16#34b# => "0010011110000000000000101100000001101101100000010000000",
16#34d# => "1000000011000111101010000000000101100100000000001010000",
16#348# => "0010011010000011101000101111000100101101010000000000000",
16#3fe# => "1010001100001000100010000000000100100100000000011010000",
16#34f# => "0010011100000000110000000000000001000000000000000000000",
16#349# => "0010011100001011100000101111000100101101010000000000000",
16#344# => "1010001110001001000000000111011000100100001000001010000",
16#3ff# => "1010001010001000100010000000000100100100000000011010000",
16#34e# => "0100101010000101110000110000000001110001100001010000000",
16#3fd# => "1011101100000000100000100111000101000011101000100001000",
16#3d0# => "1010001100001001000100000111011000100100001000001010000",
16#37a# => "0110100001010100000100000011011100101100001010000110000",
16#3c6# => "1011110111111000000000110011011100000011111000100010000",
16#3c1# => "0110001001000000011001111000001010011101100000001010000",
16#3d1# => "1010001010001001000100000111011000100100001000001010000",
16#3ca# => "0110100111010100000100000011011100101100001010000110000",
16#3c4# => "0110010101111000001000110011011100000011111000100010000",
16#378# => "1110101111101100001000010011010000011001110010100000000",
16#3cb# => "1011110101011110111001101011010001011110110000000000000",
16#3c9# => "0110010010001000101000000000110001000000000000000000001",
16#3c8# => "0110010100000000111001111100000110011101100000000000000",
16#1f5# => "0110010000000000001010110011001110110001101010010000000",
16#104# => "0111101111000101011001111000001010011101100000001010000",
16#379# => "1110101001101100001000010011010000011001110000110000000",
16#1f7# => "1011110011011000100010110011001111110001101010010100000",
16#19c# => "0111101001000101011001111000001010011101100000001010000",
16#1f4# => "1010001010001000100000000011011000100100001000001010000",
16#1f6# => "1010001100001000100000000011011000100100001000001010000",
16#37b# => "0100000111111001001000000100000010000000000000000100100",
16#22a# => "1001100010000101010001000000000001110100000000000010000",
16#229# => "1001010110001100101000101100000000110001100001000000000",
16#227# => "1001010000000101011001011100101100011101111001100110000",
16#224# => "1001001101001000101000100010000001100101111001001000000",
16#222# => "1001001100000000011001100100101010011101100000001001000",
16#3dd# => "0001000010001000000010011100001001100001100001001001000",
16#3d9# => "0110111100000101010011011100000001100101100000000110000",
16#3d8# => "1110110011000000100000011111100001000011101000100001000",
16#3d4# => "1110110110000000010011110000000001110001100000010100000",
16#22b# => "1001100100000101010001000000000000110100000000000000000",
16#228# => "1001010000001100101000101100000000110001100011010000000",
16#223# => "1001001110000000011001000001101011011100011011101001000",
16#3dc# => "0001000100001000100010000000001001100000011011011001000",
16#22d# => "0011001100001000001000110000000000110001100010000000000",
16#266# => "0001011000011000110001000000000001110100000000001000000",
16#225# => "0011001110001000000100101100000001110001100000001010000",
16#22f# => "0011010110001101101000000000000000111000000000000110000",
16#268# => "0011001110001000101000110000000000110001100010001010000",
16#234# => "0011010110011000010001110100000000011101100000000000000",
16#232# => "0001101111001011000100000000000001111000000100000000000",
16#230# => "1001100000001000000000000000000000101000011011101001000",
16#267# => "1001100110000101010001111000000000110101100000000000000",
16#235# => "0011010000011000010001110100000000011101100000000000000",
16#231# => "1001100110001000000000000000000001101000011001101001000",
16#23b# => "1100111011111100000100000000000000000000000000000111000",
16#236# => "0001110001110111000100000000000000111100000100000000000",
16#238# => "1101000011111100000100000000000000000000000001000000000",
16#237# => "0001110111110111000100000000000001111100000100001011000",
16#29b# => "1100111011111100000100111100000001111001001000000111000",
16#292# => "0100101110001000000100111000000000011111100000001011000",
16#28d# => "1100100101110000000100111111111100111111001000000000000",
16#29a# => "0001110100001000000100111100000000111001001000000000000",
16#28f# => "1100100110000000000100111111111100111111001000000000000",
16#28b# => "0100011001100000100000101000000001101010100001100000000",
16#287# => "1100010100111000100100110100000001011100100011011000000",
16#298# => "1101000011111100000100111100000001111001001001000000000",
16#296# => "0100110101110111000100110100000001110110110000000000000",
16#290# => "0100101000001000000100111000000001011111100000000000000",
16#233# => "1100100000000000000100111100000001111111000000000000000",
16#289# => "1001100010001000100000101000000001101010100000000000000",
16#28a# => "1100010010111000100100110100000001011100100001001000000",
16#299# => "0001110100000000100100111100000000111001001000000000000",
16#297# => "0100110011110111000100110100000000110110110000001011000",
16#286# => "0100101011001011000100111000000001011111100000000000000",
16#23c# => "1100001000001000000000000000000000101000011011101001000",
16#28c# => "1001111010000101010001111100000000111111000001000000000",
16#22c# => "0100011110111000000000110000000001110001100011001010000",
16#288# => "0001011100011000000100110100000001011111001000000000000",
16#294# => "0111000010001000100100110100000001110110110000000000000",
16#23d# => "1100001110001000000000000000000001101000011001101001000",
16#28e# => "1001111100000101010001111111111100111111001000000000000",
16#285# => "0001011010011000000100110100000001011111001000000000000",
16#2e3# => "0001101110000000000100111100000000111001001000000000000",
16#295# => "0111000100001000100100110100000001110110110000000000000",
16#24b# => "0101010000001000100000111000000001111001111101100000000",
16#24c# => "1101000010001000000000111000000000111001111001100000000",
16#2a3# => "0010011100000100111001110110101011110101111001000110000",
16#242# => "1101000101111100000000111000000000111001111001100000000",
16#2a6# => "0010000000001100111001110101101101110101111001000000000",
16#250# => "0101001001010000000000111000000000111001111001100000000",
16#239# => "1010100100000000011001110101101101110101111001000110000",
16#2ab# => "1100001011001000110001111111000101111101101101100000000",
16#248# => "0101010000001000100000111000000001111001111101100000000",
16#24d# => "0010011100000000000100111111000100111101101000000000000",
16#243# => "0010000110001000000100111111000100111101101000000000000",
16#2a4# => "0101001110001000000100111111001000111101101000000000000",
16#2a9# => "1100001101001000110001111111001001111101101101100000000",
16#249# => "0101010010000000100000111000000001111001111101100000000",
16#2a2# => "1010010011010100111001110101101101110101111001000110000",
16#247# => "1100001001001000110001111100000000111101100101100000000",
16#24a# => "1010001110001000100000111000000001111001111101100000000",
16#2a1# => "1010010010001100111001110110101001110101111001000110000",
16#245# => "1100001011001000110001111111000101111101101011100000000",
16#2a0# => "1100010101001000010001111100000001111101100001100000000",
16#244# => "1010001100001000000100111100000000111101100010000000000",
16#29c# => "1010001101010000011001110101101101110101111011010000000",
16#2a8# => "1100111011111100000100111111001101111101101011100000000",
16#240# => "0101010111010000000000111000000001111001111011100000000",
16#252# => "0010000010000100111001110101101101110101111011010000000",
16#251# => "1010100010001000000000111000000001111001111011100000000",
16#23a# => "1010100000000000111001110101101100110101111011010111000",
16#24e# => "0101010101010000100000111000000001111001111011100000000",
16#2ac# => "0010011000001100111001110101101101110101111011010000000",
16#246# => "1101011110000000000000111000000001111001111011100000000",
16#2aa# => "1100111001111100000100111111000101111101101011100000000",
16#29d# => "1010001110001000011001110110101011110101111011010000000",
16#2a5# => "1100111001111100000100111111001001111101101011100000000",
16#241# => "0101001101010000100000111000000001111001111011100000000",
16#24f# => "1010001011010000100000111000000001111001111011100000000",
16#2a7# => "1100111011111100000100111100000000111101100011100000000",
16#29f# => "1010010000001000011001110110101011110101111011010000000",
16#29e# => "1010010011010000011001110101101101110101111011010000000",
16#2c7# => "0011001010001101000100110000000000110001100010001010000",
16#2bf# => "0110001011001000100100000000000000111100000100000000000",
16#256# => "1110011001001101100000111100000001111101111001100110000",
16#2c5# => "0010101000111000011001111010101011111001111001000000000",
16#2be# => "0110001000000000000100000000000000111100000100000000000",
16#26a# => "0101111101000101101000110011010001000001101000101001000",
16#254# => "1110011111001101100000111010000000111001111010010000000",
16#2c4# => "0010101011011000011001111010101001111001111001000000000",
16#2bc# => "0101111010000000111001000000001011011000000000000000000",
16#26b# => "0011010010001000000100000000000001000000000010000001000",
16#264# => "1101011010000101000010110000110010110001100010000000000",
16#2cd# => "0011001010000000011001110000111000100010100000010001000",
16#2bd# => "0000001100000000100010011100000100111001100000000000000",
16#2c0# => "0101111100000000111001000000001011011000000000000000000",
16#2c6# => "0110001000000101100100110100000001111010110000000000000",
16#2c9# => "0110001100001000000100111100000000111111001000000000000",
16#2c2# => "0110010110000000100100111000000001011111100000000000000",
16#22e# => "1110000101000101101000110011010001000001101000101001000",
16#2cb# => "0100011010111000000100110000000001110001100011001010000",
16#2c3# => "0110010001001000100100111000000001011111100000000000000",
16#2b0# => "1101011010001000100000000000000000100000011101101101000",
16#2af# => "0101100001011101110011110000000000110001100010000000000",
16#3db# => "1101011010001101000110110011001001110001101001000110000",
16#2b1# => "1101011100001000100000000000000001100100011101101011000",
16#2ae# => "0101100110000000010011110000000000110001100011000111000",
16#2b5# => "1101011010001000101000111000000001111001100010000000000",
16#2b4# => "1101101100000000101101000000000001011100011101100000000",
16#2b3# => "1101101110000000000000101100000000111001000000011100000",
16#2ba# => "1101110010000000001000111000000001111001100010000000000",
16#2b9# => "1101110010001011101101100000000001000001100000001001000",
16#2ad# => "1101110010000000100000111011001101000001101000100000000",
16#2b8# => "1101011000000000110101101100000001101101100010000000000",
16#2b7# => "1101110000000000001000000000000000111000000010001000000",
16#2b6# => "1101101110001000101101000000000001011100011101101010000",
16#2b2# => "1101101000001000000000101111000101101101110000110000000",
16#2bb# => "0001000100001000001000101111010001101101101000000000000",
16#25c# => "0001000100001000000000011100000001100101100000000000000",
16#25b# => "1010111010000000010001000000000000101100000010000010000",
16#25a# => "0010110000001000100000011100000000100001100000001001000",
16#257# => "0010110110001000010001110000000000110001100010001010000",
16#259# => "0010101001011000101000110000000001110001100010001000000",
16#258# => "0010110010000000110001111000000000011101100000000000000",
16#253# => "0010110000000000001000110011110001110001101010001010000",
16#2cc# => "1010100100001000111001110000110011011101000100010000000",
16#255# => "0010110000000000110001111100000001011101100000001011000",
16#2d0# => "0110010010000000000000110000000001110001100010001101000",
16#25e# => "0110100111011101100100011110000000011101111001100000000",
16#2d7# => "1010111100001000010001101100000001101101100010000000000",
16#2d6# => "1110101110001000100000011100000000100001100000000000000",
16#2c8# => "1110101010001000010101000000000001000000000000000000000",
16#2d1# => "0110010100000000000000110011110000110001101010001011000",
16#2d5# => "1110101110001000010101011100000001100100100010000000000",
16#260# => "1110101100000000100000011100000000110001000001011010000",
16#2ce# => "1011000010000000011001000000110011101100000010000110000",
16#2ca# => "0110100000001000010001111001000000011101111001101100000",
16#2d3# => "0110010110111000000000110000000001110001100010000111000",
16#25d# => "0110100010001000010001111101000000011101111001100000000",
16#2d2# => "1010111100011000101000110000000000110001100010000000000",
16#25f# => "0101111100000000111001000000001011011000000000000000000",
16#041# => "1010010010000000110011101111000101101101110000000000000",
16#3e1# => "1010001110001001000000000100000000100100000000010000000",
16#043# => "0111000000001001001101001111010010111000001010000000000",
16#057# => "0010000001011000101000101111000101111001010010011011000",
16#054# => "0010101100001000111001000000110101011100011101100000000",
16#049# => "0010101001011000000000110000000000110001100010000000000",
16#03e# => "1010010100000000110011000000000000100100011101100000000",
16#3e9# => "1001111000001000000010110000000010110001100010000110000",
16#3e4# => "1111010110000011110011011100000001100001100001000000000",
16#3e3# => "1111001001011000000000011111100001000001110000101001000",
16#3d5# => "0111000001000000110011110011001100110001101000001010000",
16#055# => "0010101110001000111001101100111000011101100000000000000",
16#03f# => "0010101110000000101000000010000000110000011101100000000",
16#056# => "1001111010001000111001000000110010011100011101101000000",
16#3e8# => "1001111110001000000010110000000010110001100011000111000",
16#3ea# => "0111011100000000110101000000000001000000000000000000000",
16#3e5# => "1111010000001101001000111000000001111001100010000000000",
16#3da# => "1111001100000000101101000000000001011100011101100000000",
16#3ed# => "1110110010001000000000101100000000101101100010000001000",
16#3e6# => "0111011000111011110101100100000001110101100001000000000",
16#3e7# => "0010110110000000100010000000000010100000011101101101000",
16#3eb# => "1111001010001000110101101111110001101101001010000000000",
16#3ef# => "0111011100000000100000101011100000101001110000110110000",
16#3ee# => "1110110010001000000000101100000001101101100011000001000",
16#3ec# => "0111011100001000000000101011100001101001110000110111000",
16#058# => "1011000000001000011001100010101010100001111001000111000",
16#05a# => "0010110010000101101000101011111101101001001000001010000",
16#042# => "0010110110001000011001000000101011011100011101100000000",
16#05f# => "0010000110001000000000000000000001000000000000000000000",
16#059# => "1010111011011101110101101100000001101101100010000000000",
16#05d# => "0010110000000000100000000000000000111100011101101100000",
16#05c# => "0010110110000000100000000000000000111000011101101011000",
16#05b# => "0010110000001000011001000000101101011100011101100000000",
16#05e# => "0010110000001000100000000011011100101100001010000000000",
16#452# => "0010110110110000001000111100000001100101100000000000000",
16#446# => "0010101110000000100000011101000000111101111100000000000",
16#451# => "1010001010001000011001100101110101100101111001100000000",
16#450# => "1010100100110000101000111100000001100101100000000000000",
16#444# => "1010100101010000011001110101101011011101111100000000000",
16#062# => "1010001000000000000010011100010000100101111001101101000",
16#012# => "1011000011110000000100010011000101011001110001110000000",
16#0d1# => "0000100110001000011001100010101010100001111001010110000",
16#454# => "0010101110000000100000011101000001111101111100010000000",
16#453# => "0010101000000000011001100101110101100101111001100000000",
16#063# => "1010001110000000000010011100010001100101111001101100000",
16#013# => "1011000001110000100100010011000101011001110001110000000",
16#0d3# => "0000100100001000111001100010101010100001111001000111000",
16#0da# => "0110100100111101100000000000000000100000000000000000000",
16#060# => "1110011110000110100000101111101100000001101001110001000",
16#0d2# => "1011000111110000011001100010101011100001111001010111000",
16#0de# => "0010000110000000000110000000110101000000000000000000000",
16#0d8# => "0110100110111101100000011100000000100001100000000000000",
16#0db# => "1110110011101000010101101011111101101001001000000000000",
16#0ce# => "1110110100001110101000101100000001101101100000010000000",
16#0cd# => "1110011000001101010101100000000000011101100000000000000",
16#061# => "1110011000000110100000101111101100000001101001110001000",
16#0d0# => "1011000101110000111001100010101011100001111001000110000",
16#0cf# => "0110111011101000001000101111100000101101001000000000000",
16#065# => "1110011010000000100000011100000001101101100010000000000",
16#064# => "0011001000000000100100011100000000011101100000010001000",
16#0cc# => "0011001010000000011001101011111000101001001000010000000",
16#45c# => "0110100100000101101010101000000011101001100010001011000",
16#459# => "1010111100111100111001110001101101011101111100000000000",
16#4ca# => "0010101100001000111001111001101100111101111100000000000",
16#45d# => "0110100010110101101010101000000010101001100010000000000",
16#45b# => "1010111010111100111001110001101100011101111100010000000",
16#457# => "0010110010110000100000011100000001100101111001100000000",
16#4c8# => "0010101010001110111001011101101101111001111100000000000",
16#458# => "0110010111010000000000100101000001100101111001100000000",
16#45e# => "0110100010110101101010101000000010101001100010000000000",
16#4c9# => "0010101100001110111001011101101100111001111100010000000",
16#45a# => "0110010101010000100000100101000001100101111001100000000",
16#455# => "0010110000110000011001111000110011100101100000000000000",
16#45f# => "0110100100000101101010101000000011101001100010001011000",
16#4cd# => "1010111110111100110101110001000001011101111100000000000",
16#456# => "0110100000110000000000000011010001101100001010000100000",
16#4cb# => "0010101010001000111001111001101101111101111100010000000",
16#4cf# => "1010111000111100110101110001000000011101111100010000000",
16#4d0# => "1110101110000000110101011100000001110001100000001010000",
16#4cc# => "1110101000001000010101110001000001011101111100000000000",
16#4d5# => "1110011011011101000000011100000001100101111001100000000",
16#4d2# => "1110101000000000110101011100000000110001100000001011000",
16#4d4# => "0110100001011000000000101111011100000001101000100001000",
16#4d1# => "1110101000000000010101101111100001101101110000001010000",
16#4d6# => "0110100010110000101000101111100000101101110010000000000",
16#4ce# => "1110101110001000010101110001000000011101111100010000000",
16#4d3# => "1110101110000000010101101111100000101101110000001011000",
16#0d4# => "0110001110001000101000110000000000110001100000010000000",
16#07a# => "1110101100000101010001000000000000000000000000001011000",
16#0c5# => "1011110010001000000000101111001100000001101000100001000",
16#0c7# => "0110001000000000110101101100000001101101100000010000000",
16#06f# => "0110001110001000100000011100000000110001000000000000000",
16#0c4# => "1011011100001011111001000000111001000000000000000000000",
16#0dd# => "0110001111011000000000011111100001000001110000100000000",
16#0dc# => "0110111101100000110101110000000000100101100001000000000",
16#0d5# => "1111100100111101101000110011000100101101110010011101000",
16#06e# => "0110001100001100100000011100000000110001000000000000000",
16#0c6# => "1010001010001001000100000111100100100100001000001010000",
16#06a# => "0110001011011000000000100000000001000001111010100000000",
16#0d9# => "0011010000011000000100000000000001011100011011100000000",
16#0d7# => "1110110010000000110001000011100001100000010000000000000",
16#068# => "1110101000001000101000110000000000110001100010000000000",
16#0d6# => "0011010000000000010001000010000001011100011011010000000",
16#0df# => "1110101100001000000000000011010001110000001010000000000",
16#0f6# => "1000000010001001000100000100000001000000000000000000000",
16#0c1# => "0111101101011101101000101100000001101101100010000000000",
16#0eb# => "1110000010000000110101000000000001011100011101100000000",
16#073# => "1111010000001000100000010011100101011001110001110000000",
16#0f2# => "0011100001001000111001000000101010000000000001000110000",
16#0f7# => "1111010000001000100100111100000000011101100000001010000",
16#071# => "1111010011011000100000000000000001000000000000000000000",
16#0f1# => "0011100001001000111001000000101011000000000001000111000",
16#0f5# => "1111010010001000100100111000000000011101100000001100000",
16#0f4# => "0011100000000000111001000000101100000000000000001011000",
16#023# => "0011100000000000100100110100000000011101111101001010000",
16#0f0# => "0001000010001000111001000000101011000000000000000000000",
16#46a# => "1111100000001000000010000000000010000000000000001011000",
16#469# => "0011010100001000000100100100000000011101111101101101000",
16#468# => "0011010110000000111001000000101101000000000000000000000",
16#467# => "0011010010000000000000011110000001111001111101100000000",
16#465# => "0011001000001000111001111000110010100001100000000000000",
16#006# => "0011001110000000100010011110010000111101111101100000000",
16#0e9# => "0000001000001000011001111100110100100001100000000000000",
16#0f3# => "0001000010001000111001000000101011000000000000000000000",
16#400# => "1010001100001001000100000111010100100100001000001010000",
16#278# => "1000000100000011100110110000010001101101100000000111000",
16#317# => "1011110111111011100110101100001001000001100011111010000",
16#279# => "1000000010000000100110110000010000101101100000000110000",
16#314# => "0000001011001000110000110000000001110001100001011010000",
16#2de# => "1111111100001001000000011100100100101100011000000110001",
16#27a# => "0110111010001100001100000000000001011000000000000000000",
16#307# => "1010001000001001000000000111010100100100001000001010000",
16#315# => "0000001101001000110000110000000000110001100001011011000",
16#2df# => "1111111010001001000000011100100101101100011000000111001",
16#27b# => "0110111100001100001100000000000001000000000000001100000",
16#316# => "1010001100001000100110000000000110100100000000011010000",
16#178# => "0011100000001000000000000000000001000000000000000000000",
16#359# => "1011110110000100100110011110000100000001111011011001000",
16#352# => "0010110001111100001100100100000001100101100011000000000",
16#305# => "1010100011011100100000011100000000100001100000000000000",
16#17a# => "0111000111001100111001000000101111000000000000000110000",
16#179# => "1011110110001011100000111000000001111001100000010000000",
16#358# => "1101011100001000000100011110000001011101111000101001000",
16#353# => "1010100110001000000100110100000000110101100001100000000",
16#173# => "0011100010000000100100111100000000111101100000010000000",
16#17b# => "0011100100110000110000110000000001110001100001010000000",
16#3ae# => "1011110100001100100010111000000101111001100000010000000",
16#35a# => "1101011010001000000100011110000000011101111000111001000",
16#350# => "0010101111111100001100100100000001100101100011000110000",
16#171# => "1010100001010100100010011100001110100001100000000000000",
16#17d# => "0011100100110000110000110000000001110001100001010000000",
16#35b# => "1101011100001000000100011110000001011101111001111001000",
16#355# => "0010101010001000000100011110000000011101001000000000000",
16#351# => "1010100100000000000100110100000000110101100001100000000",
16#17c# => "1111100110001000111001000000001011011000000000000000000",
16#356# => "0011111010000100101010111000000101111001100000010000000",
16#357# => "0010101000001000000100100000000000011101001000000000000",
16#354# => "1010001100001000100010000000000100100100000000011010000",
16#413# => "1000000010001000001000111100000001111101100001100000000",
16#40f# => "0000100100001100101100111000000000111001100001010000000",
16#410# => "1000011010001011100000100100000001100101100011000000000",
16#407# => "0000100010000100010000000000000000000000000101101001000",
16#406# => "0000001100001000100100000010000000110100011001100000000",
16#403# => "0000001100001000000000101100000000110001111001000000000",
16#401# => "1000000110001000101100110100000001100001100000001000000",
16#412# => "1000000100001000101010000000001101000000000000000000000",
16#480# => "0000100010001000000100011111100000011100110000000000000",
16#40e# => "1010001010001001000100000111010100100100001000001010000",
16#411# => "1000011001001000000000011100000001000001100000000000000",
16#402# => "1000000010001000101100000000000001000000000000000000000",
16#481# => "1000000000001000000000111100000001111101100001100000000",
16#415# => "0100000010000100111001111000101110111001100001010000000",
16#418# => "0000111101011101101000101100000001101101100010000000000",
16#41f# => "1000110010000000010101111000000000011101100000001100000",
16#417# => "0000111000001000101000000000000000000000000000001101000",
16#416# => "1000101110001000110101101111000100101101110010011011000",
16#414# => "1000101000001000000100000011001001101100011000010000000",
16#40c# => "1000101100000011100100100100000001100101100011000000000",
16#41e# => "1000110000000000010101111100000000011101100000001010000",
16#482# => "0000100100001000000100011111001000011100110000000000000",
16#41c# => "1000110110000000010101000000000001011100000000001101000",
16#483# => "0000100010001000000100011111010000011100110000000000000",
16#41d# => "0100000100001100111001000000101111000000000000000000000",
16#420# => "1010001110001000100110000000000100100100000000011010000",
16#42a# => "1000000110001000101010000000000101000000000000000000000",
16#437# => "1001010011010101000100101100000001011111001000000000000",
16#436# => "0001101000001000101100011100000000101101100000000000000",
16#421# => "0001101000001000000100011100000001100010100000001101000",
16#35e# => "0001000001111100000010100100010001000001100000000011000",
16#37c# => "1010111100001000010000110000000001110001100011000000000",
16#42b# => "1000000000001000101010000000000101000000000000000000000",
16#438# => "1001010011010101001100000000000000100000000000000000000",
16#422# => "0001110100000000000100011100000001011111100000001100000",
16#428# => "1001100100000100101000111000000000111001100011000000000",
16#424# => "1001010101010101001100000011010101100000010000000000000",
16#423# => "1001001010001000000100011100100101011111100000001100001",
16#41b# => "1100001000110000100100100000000001011100100000001100000",
16#44b# => "1000110100001101100100111000000001111001100010000000000",
16#429# => "1010010010001000101000100111000101100101110010010010000",
16#426# => "1001010011010101001100000011111101100000010000000000000",
16#41a# => "1100001110110000100100100000000001011101000000000000000",
16#487# => "1001010101010101001100110000000001110001100011000000000",
16#485# => "1100001110001000100100111100000000111101100010000000000",
16#439# => "1100001100001000100100101100000000100010100000000000000",
16#42d# => "0001110100000000100100101110000001011111001000000000000",
16#484# => "0001011000000000000000110100000001110101100010000000000",
16#42c# => "1100001010001000010000000000000001000000000000000000000",
16#435# => "1100001100001000100100101100000001011100100000000000000",
16#43b# => "1100001110001000100100011110000001011111001000000000000",
16#486# => "0001110110001000100000101100000001100000100000000000000",
16#434# => "1100001110110000010000100100000001100101100010000001000",
16#42e# => "0001101000000101000100110000000000110001100010000000000",
16#433# => "0001011101111100000000011100000000101101100000000000000",
16#431# => "1001100110001100110000100111000101100101111010010011000",
16#488# => "1100001100110000100100101110000001011110110000000000000",
16#43a# => "1100010100000000000100111000000001111001100010000000000",
16#425# => "0001110110001000001000100111000101100101110010010010000",
16#42f# => "1001001111010000101100101110000000011100110000000000000",
16#432# => "1001100010001000100000111100000000111101100010000000000",
16#430# => "1001100000000000100100110100000001110101100010000000000",
16#427# => "1000000000001000101010000000000101000000000000000000000",
16#112# => "0101010000000000100100000000000101110100000000011110010",
16#1a9# => "1011110000000001011001000000010110000000000000000010000",
16#111# => "0101010100000000100100000011000110110100001000011110010",
16#079# => "0001011100000000100000011100000001100101100000001100000",
16#113# => "1011110110000001011001000000000011110100000000000010000",
16#01f# => "0001011000001000100100000000111001000000000000000000001",
16#017# => "0000111010001000100100000000000001100101100011111100100",
16#110# => "1000101110001011100110100010000010011101111000000000000",
16#01e# => "1001010110000000000100101111110100101101101010000000000",
16#026# => "0000111100001000000100000011011000101100010000000001000",
16#02c# => "1001001000001000000100100000000000100001111000000000000",
16#016# => "0001011100000000000100011100000000100001111000000000000",
16#02e# => "1001010010111100100000101111010101100010101001110001000",
16#01d# => "0001011010001000000100011110000001011101111011100000000",
16#028# => "0000111110000101010100101100000001101101100010000000000",
16#01c# => "1001010000111000100000000000111101000000000000000000001",
16#02a# => "0000111000000101010100101100000001101101100010000000000",
16#029# => "1000000101000111100110000000000101000000000000000000000",
16#030# => "0001110110000000000100000011001100101100011000000000000",
16#031# => "1001100000000000001000110000101101110001100000000000001",
16#039# => "1001100110000000110100001000000001011101100000000100100",
16#027# => "1011101110000000100100000011100000101100010000000001000",
16#1ba# => "1011101110000001000000000011001011101100011000010000000",
16#03b# => "1001100100001000010100110100000000011101100000001100000",
16#075# => "1011101000001000100100000000000000110100000000000000000",
16#02d# => "0001101110001000100100000011110001101100010010000001000",
16#087# => "1010100111010000001000101111100000101101101000001000000",
16#085# => "1100001000001101110100101100000001101101100010000000000",
16#084# => "1100001110000000100000111100000001111101100000000000000",
16#03a# => "1100001010000000011001111000100100111001100000000000000",
16#032# => "0001110100001101101000101100000001101101100010001100000",
16#038# => "1001100000001000010100100100000001011101100000001101000",
16#077# => "0001110110000101000100000000000001000000000000000000000",
16#037# => "1011101101010000100100101111010001101101101010010000000",
16#02f# => "0001101100001000100100000011111001101100010010000100000",
16#086# => "1001100000001000101000101000000000101001100000001101000",
16#033# => "1100001010000000011001100000100010100001100000000000000",
16#147# => "0001101000001001000100000011110111101100010010000100000",
16#08a# => "0100011000000000010101111100000000011101100000000000000",
16#1f0# => "0011010000001000010101111000000000011101100000000000000",
16#1e7# => "1111100100000101100000011100000000101011100000000000000",
16#16b# => "1111001010001000100100011100001001011100100000000000001",
16#08b# => "0100011111011000010100111100000000011101100000000000000",
16#16a# => "1100010100001101101010101100000011101101100010000000000",
16#1f1# => "0011010010001000010100111000000000011101100000000000000",
16#381# => "1111100010000101100010011100000101100011100000000000000",
16#159# => "0100000001000001011001001100101110100100000000000100000",
16#021# => "0010110010000000100010010000000100011001110000110000000",
16#050# => "0001000010000000111001010011010000011001110010100000000",
16#383# => "1101011000001000100010011100000101100011100000000000000",
16#052# => "0100000000000001011001001101101111110000011000000000000",
16#08f# => "0100101100000000010100000000000001000000000000001010000",
16#08d# => "0100011010001000100000000000000001000000000000000000000",
16#089# => "0100011100000000111001000000000001000000000000000000000",
16#08e# => "1100010110000000101000101100000001101101100010000000000",
16#094# => "0100110101100110001000101010000001101001001000000000000",
16#091# => "0100101100000000010100000000000001011100000000010000000",
16#090# => "0100101110000000010101000000000001011100000000010000000",
16#08c# => "1100100000001101101000101100001101101101100010000000001",
16#093# => "0100101010000000010100000000000000011100000000000000000",
16#092# => "0100101000000000010101000000000000011100000000000000000",
16#036# => "0001101010000000001000110011000101100101101000100000000",
16#018# => "0001101011001000010101110100000001111101100000000000000",
16#034# => "1000000000000111101010110000000100111001100000000000000",
16#01a# => "0001101100000000010101111000000001110001100000000000000",
16#098# => "1100111001110111000100100011010001100010110000000000000",
16#03c# => "1011101110001000101010110011001111110001101010000000000",
16#019# => "1001111100000000010100101111010000110001110000000000000",
16#095# => "1000110111010101100100100011001101011101110000000000000",
16#09c# => "0100101111111000100100101100000001101101100010000000000",
16#099# => "1100111111110111000100100011100001100010110000000000000",
16#097# => "1000110101010101100100100011001001011101110000000000000",
16#09d# => "0100101100001000000100100011000101011101110000000000000",
16#09a# => "1100111111110111000100100011100001100010110000000000000",
16#09f# => "1100001110001000101010101011010110101001101000000000000",
16#01b# => "1100111110001000110100000011000100101000010000110000000",
16#096# => "1000110111010101100100101100000001101101100010000000000",
16#09e# => "0100101000001000000100100000000000011101100000000000000",
16#09b# => "1100111101110111000100100011110001100010110000000000000",
16#3b1# => "1010001110001001000000000100000000100100000000011010000",
16#324# => "0101100010000100011001000000100101000000000000000000000",
16#3b6# => "1010001100001001000100000111010100100100001000001010000",
16#3b0# => "1101101101001000000000011111000101000001101000101100000",
16#326# => "0101100000000000011001010100100100100001100000000000000",
16#3b8# => "1010001110001001000100000111001000100100001000001010000",
16#3b4# => "1101110111111011100100110011011101000011110000100010000",
16#325# => "0101100000000000011001000000100101000000000000000000000",
16#3bc# => "1010001000001001000000000111011000100100001000001010000",
16#3ba# => "1010001000001001000100000111001000100100001000001010000",
16#3bd# => "1000000110000000000000100000000101010101100000000000001",
16#3bb# => "0101111111010100010000010111010001010101110010101101000",
16#3bf# => "1000000000000000000000100000000101010101100000000000001",
16#3de# => "1101101110000000100000110000001101110001100000011110000",
16#3b9# => "0110111000001111010000000000000001000000000000001100000",
16#03d# => "1101000100001000100100011100000000001101000000000000000",
16#0a1# => "1001111100000000101000011111001001000001111000100001000",
16#0a2# => "1101000100000000111001011101100100000011111000100010000",
16#35c# => "1101000110001000000010000000000010000000000111110000000",
16#3b7# => "1010111110000000010000110011001100110001101000001010000",
16#3b3# => "1101101100001000101000000011010000100100010001001000000",
16#3b5# => "0101100000001101111001101000100010100001100000000110000",
16#3be# => "1101101110000000100000110000001101110001100000011110000",
16#377# => "0101111010001000010000000000000001000000000000000000000",
16#3b2# => "1000000011000111101010000000000101100100000000001010000",
16#0a6# => "1000000111000111100010000000000101100100000000001010000",
16#0a8# => "0101001000001101100100100011100000011100110000000000000",
16#070# => "1010001000001000100000011100000000100001100000001001000",
16#048# => "0011100011010000010000110011001000110001101000000000000",
16#0a7# => "1010010101011100101000001000000001000001100011000000100",
16#0a9# => "0101001110001101100100100011010000011100110000000000000",
16#0a4# => "0101010001111100011001011100101110100001100000000110000",
16#053# => "0101001010000000000000011110000000101010110000000000000",
16#0a3# => "1010100110001000110000110000000000110001100000010000000",
16#072# => "1010001110001000100000011100000001100001100001001001000",
16#0aa# => "0101001110001101100100100011001000011100110000000000000",
16#051# => "1010100000001000110101101000000000100001100000001100000",
16#0ab# => "0101001000001101100100100011000100011100110000000000000",
16#046# => "0101001100001000111001100000000001011101100000001011000",
16#044# => "1010001010001000000000011100000000111001100000000000000",
16#047# => "1010001010000011110000110000000000110001100010000000000",
16#04d# => "1000000110000111100010011100000101111101100000000000000",
16#04a# => "0010011101000101010000111011000101100101101000101001000",
16#045# => "1010010100001100100000011100000000111001100000000000000",
16#04f# => "1111100100001000000010011100000101111101100000001100000",
16#1f2# => "0011010010000000111001010011010000011001110010100000000",
16#04e# => "1111100010001000000010011100000101111101100000000000000",
16#04c# => "1001010000001000100000011100000000111101100000000111000",
16#0f9# => "0101100110001000100000011100000001111101100000000000000",
16#04b# => "0111110110000000110000010111010000010101110000111100000",
16#0fa# => "1001001010000011100100000000000000000000000111110000000",
16#0ef# => "0111110100001101100000011111001001000001101000100000000",
16#0c0# => "0111011110001000111001111001100101100101101000101001000",
16#0a0# => "1110000011010000000000010011001110011000111000101110000",
16#0a5# => "1101101010001000011001000011100011100100010000010000000",
16#0ad# => "0101001100000000100000011100000001100001100000000010000",
16#088# => "1101011010000000111001000100101111111101100000000000100",
16#015# => "1100010000000000001000000000010000111000011000000000001",
16#001# => "1000101000000000111001000000010000011100000000001100000",
16#00a# => "1101011010000000111001000000101110000000000000001101000",
16#0fb# => "0111110000000000000100101110000001000001111000000000000",
16#0ed# => "1110000110000000001000000000101111000000000000000000000",
16#0c2# => "0111011100000000111001100001101110011100110000000000000",
16#0b6# => "1101000100000000000100011100000000101101100000001010000",
16#0f8# => "1101011000000000000100000000000000000010000000000000000",
16#005# => "1101011010111000000100000000000001000000000000000000000",
16#0bc# => "0000001100000000100100010100000000010101100000001000000",
16#0ac# => "1000000110000000000110000000000101000000000000000000000",
16#0ff# => "1101011010111000000100111010000000000010011000000000000",
16#078# => "1111111110001000100100010100000000010101100000001101000",
16#0bd# => "1011110110000000000100111100000000100001100000001010000",
16#024# => "0101111110000000100100011100000001001101000000000111000",
16#0af# => "1000000110000111100110000000000101000000000000000000000",
16#025# => "0101111000000000100100011100000000001101000000000000000",
16#10d# => "1001010110001000100010011100000011101011100000000111000",
16#0ae# => "1101011100001111100100111010000001000001100110110000000",
16#02b# => "1101011010001000000100111100000000100001100000000000000",
16#0e4# => "1111001010000000100100000000000000100000000000000000000",
16#0e5# => "0011111000000000000100100011001001000001101000000001000",
16#074# => "1111001010000011100100000000010001100000011000001011001",
16#080# => "1011101000000000000100000111111101000001111001110010100",
16#06d# => "0101111000001000100100111100000001000001111010011001000",
16#0e2# => "1011011010000000100000011100000001110101100000001101000",
16#0bf# => "0111000101011101110101101100000001101101100000010000000",
16#07c# => "0101111000110000100100000011010000101100011000001100000",
16#0be# => "0101111011001000100100111100000001011101100011011100000",
16#06b# => "0101111000001101000100111000000001000001111010011001000",
16#0e3# => "0011010000001000100000011100000001110001100000001010000",
16#076# => "0101111100000011100100000000000000000000000000001000000",
16#00f# => "1011101110001000000000011110000000000001111001110000000",
16#069# => "1000011110001000110000000000000001000000000000000000000",
16#0e1# => "0011010010000000100000011100000000100001100000000000000",
16#007# => "0101111101010100100100111000000000011101100001000100000",
16#0e0# => "0000001000001000101000000000000001000000000000000000000",
16#0c8# => "0111011100000000000100000000100110101100000000011110000",
16#07b# => "0110010110001000111001000000110000011000000011010000000",
16#0e7# => "1011110010001000101000110011001001110010110010000000000",
16#0fe# => "1111010000000000001000101111100001101101101000000000000",
16#022# => "1111010010001000001000000000111100011000000000001110000",
16#0ca# => "0001000110001000011001000000010001010100000000000000000",
16#0cb# => "0110010001010100101000110011110001110001101000000010000",
16#0e6# => "0110010000011000101000110011000100000001010001000000000",
16#0c9# => "1111001010001101110001110000000000110001100000010000000",
16#0ee# => "0110010110000101000100010011001000011001111000010000000",
16#0e8# => "0111011110110000000100000011100101110000011000000000000",
16#0ec# => "1111111100001000010110000000000001001100000000000000000",
16#ab8# => "0111011010000000000110000000000011101100000000010000001",
16#328# => "0101111010001000010000000000000001000010000000001101000",
16#0ea# => "1001010000000000000110000000001111110000000000000000000",
16#aba# => "1000011000000000000110000011101100101000000001110011000",
16#abb# => "1101110111001000000100000000101101111000000000001000001",
16#014# => "1101110110001011100110001000101010011110100000001001100",
16#00e# => "1000101100000000001000000011100001000000101010101111000",
16#000# => "1000011110001000010110011011100001011100010000000000000",
16#0b3# => "1001001000001000100100000000000001100100000000000110000",
16#0b2# => "0101100010001000000100000000000000000010000000000000000",
16#0b1# => "0101100010001011100100010111010001010101010000111010000",
16#083# => "0101100000000011100100010111010000100001110000100000000",
16#00d# => "0100000000001011100000010111001001000001101000101100000",
16#004# => "1000011000000000111001010111010001000001101000100000000",
16#1fe# => "1110011010000000100100000000101101100100000000000000001",
16#1ff# => "1111111000001000000100010111010000010101110010100000000",
16#0bb# => "1011011110000000000100011111010001000001110000100000000",
16#0b5# => "1101110101010011100100010100000001010101100000000000000",
16#035# => "1101101010000011100000010111001001000001101000100000000",
16#020# => "0001101000000000111001010111010000000001101000100010000",
16#0b9# => "1010001000001001000100000111010000100100001000001010000",
16#0b4# => "0101010010001000000110010100100111010101100000000000000",
16#040# => "0001101000000000111001010111010000000001101000100100000",
16#18a# => "1100010010000000000100011100000000011101100001100000000",
16#16d# => "1100001011011000011001000000000000011100000000011011000",
16#120# => "1011011111001100100100000000000001101000000000000000000",
16#188# => "1010001000001000101000000011010100100100001000000000000",
16#16c# => "1100010000000000011001000000000000011100000000011011000",
16#122# => "1011011101001100100100000011010000101000010000001010000",
16#11e# => "0001000100111000000100111100000001111101100001101001000",
16#07f# => "0000111100001011100110111000000100111001100001010000000",
16#06c# => "0011111110001011100100111011000100000001101000101000000",
16#16e# => "1010001110001000100100000011010100100100001000000000000",
16#11f# => "1011011110001000000100111000000001111001100010001010000",
16#07e# => "1010001010001001000100000111010100100100001000001010000",
16#365# => "1010001110001001000100000111011100100100001000001010000",
16#81c# => "1010001110001001000100000111011100100100001000001010000",
16#829# => "0000111010001010100100000000000000011100000000000000000",
16#828# => "1001010000000000100000110000000001110001100011000000000",
16#36c# => "1001010010000000000110100000100001011101000000000000000",
16#360# => "1011000110001000000000101011001100101001110010100000000",
16#81e# => "1010001000001001000100000111011100100100001000001010000",
16#36d# => "1001010100000000000110100000100000011101000000001101000",
16#36b# => "1011011001101000101100011100000001100001000000000000000",
16#364# => "0011010001011011100100011111110101000000101010011100000",
16#362# => "0011001100000010100000011111101101000000101010010110000",
16#37e# => "1011000011111100010000100100000000101101100000000011000",
16#820# => "0001000110000000100100110100000001110101100010000000000",
16#36f# => "1011011110001000000000010011100000011001110001111101000",
16#36a# => "1011011111101011101100011100000001100001000000000000000",
16#361# => "0011001100000010100000011111101100000000101010010111000",
16#821# => "1001001100001101100100011110100101100011010111101001001",
16#81f# => "0001000110000100100100010011100000000001110001001011000",
16#36e# => "0011001100000010100000011111101101000000101010011010000",
16#363# => "1011000010000000100000101011000100101001101010100000000",
16#367# => "0011001100001000000100010011100000011001110001111101000",
16#369# => "0011001110001000100100011110000001011110110000000000000",
16#366# => "0000111011110010100110110000100001110001100011000000000",
16#368# => "0011001000001011100100011110000001011110110000000000000",
16#800# => "1010001000001001000100000111011100100100001000001010000",
16#726# => "1000000110000010100010011100100000100001100000000000000",
16#720# => "1001001110110000010000101111000100101101111010010011000",
16#824# => "0001000000001100001100100011101000011101001000000000000",
16#728# => "1010001100001001000000000111011100100100001000001010000",
16#804# => "1001010110110000100110100000011100011101100000001001000",
16#801# => "0000001011101100001100110000000000110001100010000000000",
16#724# => "1001001000001000000000111100000000111101100010000000000",
16#822# => "0001000101010101001010111000011100111001100010000100000",
16#825# => "0001000010001100001100100011101100011101001000000000000",
16#72a# => "1010001010001001000000000111011100100100001000001010000",
16#806# => "1001010000110010100110011110011100011101111111101001000",
16#80e# => "0000001011101100001100101111000100101101110010010010000",
16#721# => "1000011000110000000110000000100001100000000000000001000",
16#823# => "0001000111010101000010111000011100111001100010000100000",
16#826# => "0001000110001100001100100011110000011101001000000000000",
16#729# => "1001010110001000100000110100000001110101100010000000000",
16#807# => "1001010110110010100110011110011101000001111111101001000",
16#80c# => "1000011100001000000100111100000000111101100010000000000",
16#827# => "0001000100001100001100100011110100011101001000000000000",
16#72b# => "0001000001010101000000111000000000111001100010000100000",
16#723# => "0011100110111100100100111000000001111001100000010000000",
16#730# => "1010001000001001000100000111011100100100001000001010000",
16#72c# => "1001111110000000000100000000000001000000011111101001000",
16#722# => "0010000100000000110000110000000000110001100010000000000",
16#736# => "0001101100000000000100100000000001000001100000000000000",
16#732# => "1010001110001001000100000111011100100100001000001010000",
16#72d# => "1001111000000000000100000000000000000000000011010000000",
16#741# => "1001100000110010100000101100000000101101100010000001000",
16#737# => "0001101010000000000100100000000001000001100000000000000",
16#738# => "0001000010001101000100000011111100000000011101011010000",
16#735# => "0001101100000000000100100000000000000001100000000010000",
16#73c# => "0001110100000011100100000000000001000000000000000000000",
16#72e# => "1001111100001000000100000000000000100000011111101001000",
16#731# => "0001011110111100100100110100000001110101100010000000000",
16#739# => "0001000100001101000100000000000001000000000000000000000",
16#734# => "0001110010000011100100000000000001000000000000000000000",
16#73e# => "0001101011010100100100100011100101000001111010010000000",
16#72f# => "1001111111001000000100000000000000100000011111101001000",
16#733# => "0001011100111100100100000000000001000000000000000000000",
16#782# => "1011101100000000100100011111001000011100110000000000000",
16#770# => "0100000011001101111001100100101110100111100000000000000",
16#783# => "1011101010000000100100011111010000011100110000000000000",
16#773# => "0100000011001101111001100100101110100111100000000000000",
16#775# => "1001111010001000100000000000000001000000000000000000000",
16#780# => "1011101010000000100100011111100000011100110000000000000",
16#774# => "1011101100001100000000111001000000111001101000000111000",
16#781# => "1011101100000100000100011111100000011100110000000000000",
16#777# => "0011100000001000100100010011000101011001101001110000000",
16#772# => "1011101000000000000100100100000000100111100000000000000",
16#784# => "1010001000001001000000000111101000100100001000001010000",
16#7ed# => "0011100100001000100000000000000000000000000010001001000",
16#785# => "0000001010000000100010011100000100111001100000000000000",
16#73f# => "1100001100000011111001000000001011011000000000000000000",
16#7ef# => "1001111010001000100000011111010001000001101000100000000",
16#7ec# => "0111011110001000100100011111000100011100110000000000000",
16#771# => "0111011100000100011001000000101111000000000000000000000",
16#77a# => "1011101110001000000000111100000000111101100000010000000",
16#7ee# => "0011111000000101001100100000000000011101001000000000000",
16#7e7# => "0111011100001000000100011111000101011100101001110000000",
16#778# => "1111001100001000100000000000000001100000010111010000000",
16#776# => "1011110010110000001100100100000000000001100000000001000",
16#77d# => "0011111001011000101000010011000101011001101001110000000",
16#815# => "1000110010001000100000111100000000111101100010000000000",
16#81b# => "1000101100001000101100000000000001000000000000000000000",
16#77c# => "1000110110001000001010111000100001111001100010000000000",
16#817# => "0011111100000101000100000000011100011100011111100000000",
16#81a# => "1000101110110000101100100100000001100101100010000001000",
16#3e2# => "0011111010000000100000101011100000101001101000110000000",
16#3e0# => "0011001100000010100000011111101101000000101010010110000",
16#37f# => "0111000101111000010000101011100000101001101010100000000",
16#79d# => "1010001010001001001000000111011000100100001000001010000",
16#792# => "0100101110001000000100101011100001101001110010101011000",
16#793# => "1100100000001000001000101111111101101101110000000000000",
16#78d# => "1010001100001001000100000111011000100100001000001010000",
16#78a# => "1100010010001000100100110100000001110101100010000000000",
16#79c# => "1010100000111000001000100101000001100010101010010000000",
16#796# => "1100111100000100110101100000000000011110100000001001000",
16#791# => "0100101111011000001000101100000001101101100010000000000",
16#78c# => "1100100111010000110101100000000001011101000000000000000",
16#78b# => "0100011100000100100100100101000001000011010011010000000",
16#81d# => "1100010100001100100110100111011100101100101011000000000",
16#78e# => "1010001100001001000000000111011100100100001000001010000",
16#790# => "0100101000000000001000101111111001101101101000000000000",
16#797# => "1100100110000101010101011110000001011111001000001001000",
16#78f# => "0100101010001000101000101111100101000001111001110001000",
16#79a# => "0100011000001010110101101111111100101101110000010000000",
16#795# => "0100110000110000000000100000000001100010110000000000000",
16#794# => "0100101010000000110000110000000001110001100010001011000",
16#798# => "0100110110001000000100110100000001110101100010000000000",
16#751# => "1011000010001000000100101110000001101101001001000000000",
16#753# => "1111001000001000000100100111100000101111011001000111000",
16#755# => "1010100001011000100100111100000000111101100011100000000",
16#752# => "0010101010000100000100111010000001111001111011010000000",
16#756# => "1010001000001001000100000111011100100100001000001010000",
16#75c# => "0010101100001011100100111000000001111001100010000000000",
16#75b# => "1010111111010000000000011100000001000001100000000000000",
16#757# => "0010110110110000101100100011000100100001110010010010000",
16#758# => "0010110010001000000100111100000000111101100010000000000",
16#754# => "0010110110110000000000100110000000100011001000000010000",
16#750# => "1010100000001000000100101011010000101001110010100000000",
16#760# => "1010001000001001000100000111011100100100001000001010000",
16#75e# => "1011000010000011100100111001000000110001101001010000000",
16#759# => "0010110000001000000000111100000000111101100010000000000",
16#75a# => "0010110100001000101100101101000001101101101000110000000",
16#761# => "0100110010000000100100111100000000110101100001100110000",
16#799# => "1101000000000000010000101110000001101111001000000000000",
16#7a6# => "0100110000001000101000110000000000110001100000010000000",
16#7a5# => "0101001100001101010000000000000000011100000000000000000",
16#79e# => "0101001110000010101000111100000001111101100001100000000",
16#7a3# => "1100111100001101001100111000000000111001100001010000000",
16#7a0# => "1101000101001000100000100000000000100001100010000001000",
16#79b# => "1101000110110000010000000000000001000000000000000000000",
16#7a7# => "1101011011010000001000100011010101000001110010011000000",
16#7a4# => "1010001110001001000100000111011100100100001000001010000",
16#7a8# => "0101001010000010101000011100000000100001100000000000000",
16#7a9# => "0101010000000000001100011100000000011101000000000010000",
16#79f# => "0101010000000000101000111000000001111001100010000000000",
16#7a1# => "1101000110001000100100000000000000011100000000000000000",
16#7a2# => "0100110110001000100000110100000001110101100000010000000",
16#7b8# => "1010001100001001000000000111011100100100001000001010000",
16#7c4# => "1110011011010000000000111001000001111001101001010000000",
16#7bc# => "1101101110001000010001110000000000110001100010000000000",
16#7ba# => "1010001010001001000000000111011100100100001000001010000",
16#7c6# => "0110001000000000000000011111100100000001010010010010000",
16#7c0# => "0110001100111100000100011111100101011101110111100011000",
16#7be# => "1101101000001000010001110000000000110001100010000000000",
16#7b9# => "1101110010001000100000111100000000111101100010000000000",
16#7aa# => "1101110000110010100100011110000001011101111111101000000",
16#7b7# => "0101010100001000001100111000000001111001100010000000000",
16#7b6# => "1101101011100000100000011100000000100001100000000000000",
16#7b0# => "1101101110111000010001110000000000110001100011000100000",
16#7c5# => "0011001000001101000000111001000001111001101001010000000",
16#7c1# => "0110001010111100000100011111100101011101110111100011000",
16#7bf# => "1110000011011100101100101100000001000000100010001001000",
16#7bb# => "0101111101101101000000110011100001000001111001110001000",
16#7b5# => "1101101110001000100100000000000000000000000000000001000",
16#7b4# => "1101101101100000100000011100000001100001100001000000000",
16#7b1# => "0101100000000000000100111100000000111101100000010000000",
16#7af# => "1101011000000000101000011111100101000001111010010011000",
16#7c7# => "0011001110001101000000111001000001111001101001010000000",
16#7ad# => "0110010111010101001000111001000001111001101001010000000",
16#7b2# => "1101011100111000101100011110000000011101001000000011000",
16#7c2# => "0101100110001100000000011111100101100001101110000000000",
16#7ab# => "1011000010001100101000111001000001111001101001010000000",
16#7b3# => "0101010010001000101100011110000000011101001000000000000",
16#7c3# => "0101100000001100000000011111100100100001101110010000000",
16#7cc# => "0101100100000100100100101111111100110010110000000000000",
16#7d0# => "0111000010111000000100100100000000100010100000000110000",
16#7ce# => "0110100111001000000100111001000000111001101010000000000",
16#7d2# => "0110100000000000100100111000000000111001100011000000000",
16#7cf# => "0110100001001000000100000000000001000000000000000000000",
16#7cb# => "0110100111001000000100111001000000111001101010000000000",
16#7cd# => "0110111110110000000100000000000001000000000000000000000",
16#7c9# => "1110011000000000100100011111010101000001010010011010000",
16#7c8# => "0101100110000100100100101111111000110010110000000000000",
16#7ca# => "0101100000000100100100101111111000110010110000000000000",
16#7d4# => "0110100100001000100000111100000000111101100010000000000",
16#7d1# => "1110101100111100101100101100000000101101100010001000000",
16#7dd# => "0101100000000100100100101111111000110010110000000110000",
16#7d3# => "1110101010111000101100000000000001000000000000000000000",
16#7d6# => "0110100010001000100000111100000000111101100010000000000",
16#7df# => "0101100110000100100100101111111001110010110000000111000",
16#7da# => "0110111010110000100100111001000000111001101001011011000",
16#7d5# => "1110110110000000000000011100000001000001100000000011000",
16#7dc# => "0101100010000100100100101111111100110010110000000110000",
16#7ac# => "0110111000110000000100111001000001111001101001011010000",
16#7db# => "1101011101010000000100011111010101000001010010010000000",
16#7d8# => "1110110000001101000100011111010100000011010010010000000",
16#7d7# => "1110110000000000000000011111100101000001111010010011000",
16#7de# => "0101100100000100100100101111111101110010110000000111000",
16#7ae# => "1110011010001000100100101100000001000000100010001001000",
16#7e0# => "1010111010000000100100111010000001111001111001000000000",
16#7bd# => "0111000000111100000100100100000001100010100000010000000",
16#7e1# => "1010001000001001000100000111101100100100001000001010000",
16#7e6# => "1011000010001000100100101011001001101001110010101011000",
16#7e2# => "1111001100001000000100111001000000111001101001000110000",
16#7ea# => "1111001010000000000000111100000000111101100000010000000",
16#7e8# => "1100111100000000000100011100000001011101000000001010000",
16#7e4# => "1111010000110000001100101011001000101001110000110000000",
16#7e3# => "1111001110000100100100111010000000111001111000000000000",
16#7e5# => "0101010110001000100100111010000000111001111010010110000",
16#764# => "0101100010000100100100101111111100110010110000000110000",
16#762# => "0011001010000100100100111000000000111001100001011010000",
16#765# => "0011001000000000000100111100000000111101100000010000000",
16#763# => "0101100000000100100100101111111000110010110000000000000",
16#76a# => "1000000000001001000000000100000001000000000000000000000",
16#76c# => "0011010100001100000100011111101000011101001000000000000",
16#766# => "0101100100000100100100101111111100110010110000000000000",
16#76d# => "0011010110001100000100011111101100011101001000000000000",
16#75f# => "0101100000000100100100101111111001110010110000000111000",
16#767# => "1010111111001000100100101100000000101101100010001011000",
16#76e# => "0011010010001100000100011111110000011101001000000000000",
16#769# => "1011011000001101101100000000100101000000000000000000001",
16#75d# => "0011010010000100000100111100000000111101100101100000000",
16#7d9# => "1010111010000000100100111001000000111001101011000111000",
16#76b# => "1110110010000000100000101011000100101001101010100000000",
16#76f# => "0011010000001100000100011111110100011101001000000000000",
16#768# => "1011011010001110001100000000100101000000000000000000001",
16#7fc# => "0100000101001101111001000000101110101000000000010000000",
16#7f8# => "1010010110001101101100111000000000111001100001010000000",
16#7f6# => "0111110101010101000100011111001100000000101010010100000",
16#7f4# => "0111101110001000000000011111001000000001110010010011000",
16#7fe# => "0111101010000000001100000000000001000000000000000000000",
16#832# => "1111111110110000000110111100011101111101100001100000000",
16#77b# => "1010010000001101101100111000000000111001100001010000000",
16#7f9# => "1010010000001101101100111000000000111001100001010000000",
16#7fd# => "0111101010000101100100000011010101100000010000000000000",
16#82b# => "1010010100001000100110101100011101011101100000001000000",
16#83c# => "1001010000001000101100111000000000111001100001011100000",
16#779# => "1001111010000011100110000000100001000000000000000000000",
16#7fa# => "1011110000110000100100011100000001000000100010000000000",
16#7ff# => "0111101100000101100100000011111101100000010000000000000",
16#727# => "0010011001010101101100000000000000000000000001001010000",
16#83d# => "1001001111011000100110101000011101101011000000000011000",
16#746# => "1010001110001001000100000111011100100100001000001010000",
16#73d# => "1010001110110000000100101011011001000011010001000000000",
16#740# => "1001111010000000100100101011011001000001010000000000000",
16#7f3# => "0010000000110000000000011100000000101001100000000010000",
16#725# => "1111100111000000110000110000000001110001100000011011000",
16#7fb# => "1001001111011000100100101000000000101011000000000010000",
16#742# => "0010000100000000000100110100000001110101100000010000000",
16#7f1# => "1010001110001001000000000111010100100100001000001010000",
16#74a# => "1010010010001000100100101100000000011101100000000000000",
16#83e# => "1100001110001100100010000000011101000000000000000000000",
16#74e# => "1001111000001101000110101100100000011101100000000000000",
16#74b# => "1001100000001000000010100100100000100101100010000000000",
16#786# => "1010010110001000100000111000000000111001100001010000000",
16#83f# => "1100001000001100100010000000011100000000000000001101000",
16#7eb# => "1010010100001000100100111000000000111001100001011010000",
16#74f# => "1100001110001100100100100000000001011101000000000000000",
16#744# => "0010011101010101101100101011110101000011010010010010000",
16#749# => "1001100010001000000110100100100000100101100010001100000",
16#7e9# => "1010010111010000100100111000000000111001100001011010000",
16#787# => "1111010101010000100000101011101101000011010010010010000",
16#74d# => "1100001000001100100100101010000001011110110000001001000",
16#747# => "1100010000000000010101111100000000011101100000000110000",
16#7f5# => "1100001000001100100000000000000000000000000000001101000",
16#789# => "1111111110001000101000100000100100101101100000000000001",
16#745# => "1100010110000000110101111000000001011101100000000111000",
16#788# => "1010001100111000101000101100000001101101100000010000000",
16#743# => "1100010110000000010101000000000000011100000000000000000",
16#748# => "0010000100001000100100000011000100101100011000000000000",
16#7f7# => "1010010110000000000000101100000001100001100000001101000",
16#74c# => "0111101010111000100100101010000001011110110000001001000",
16#2e6# => "1010001110001001000000000100000000100100000000011010000",
16#14a# => "1010001010001001000100000100000000100100000000011010000",
16#14b# => "1010001100001001000100000100000000100100000000011010000",
16#b1f# => "1001001111011101100100101011111101100101111001110111000",
16#b09# => "0000111001100110000100010011011101011000110001111011000",
16#b08# => "0000010111011000100100000011111101101000000011110110000",
16#b07# => "0000010010000101100100000011000000111100011001111001000",
16#b15# => "0000001110011011100100000010101100101000000111111001001",
16#b33# => "1000101100111011100000011100100001100111100001111111000",
16#b0c# => "1001100101010101000100101111111101011100000001110111010",
16#bff# => "1000011100000000010110101111111100101000000001110011000",
16#b26# => "0000111011101110100100101001000000011100011011111010000",
16#b1c# => "0000010010000000100100000000000000101010000011111100000",
16#b0b# => "0000010110000000000100000000000001000010000001110000000",
16#b05# => "1000101100000000100100000000000001110010000001110000000",
16#b17# => "1111111000001000100100000000000000101010000000000110000",
16#b32# => "1001100010001000100000000000000001000010000001110000000",
16#b0d# => "1000011010000000000000000000000001000010000001110000000",
16#b24# => "0000111101110111000100000011111100010000000001111101001",
16#b1d# => "0000010100000000100100000000000000101010000011111100000",
16#b06# => "1111111000001000100100000000000001000010000001110000000",
16#b16# => "1001100110001000100100000000000001000010000001110110000",
16#b31# => "1001100010001000100000000000000001000010000001110000000",
16#b0e# => "1000011010000000000000000000000001000010000001110000000",
16#b25# => "0000111011111100000100000011111100000000000011111011000",
16#b1e# => "0000010100000000100100000000000000101010000011111100000",
16#b14# => "1000011000000000000100000000000001000010000001110000000",
16#b30# => "1001100100001000100000000000000001000010000001110000000",
16#bfe# => "1101110110001000100100000000000001000000000000000000000",
16#b58# => "0001011111011000100100000011111101000000011001111011000",
16#b1a# => "0010110010000000000100111000000000111001100001110111000",
16#b2c# => "1000110010100000000100000011111101001000001001110001000",
16#b11# => "0001011101001000000100000011010001010000010001110010000",
16#b12# => "0000100000000000100100000011000101101000001011111000000",
16#b0f# => "0000100100001011100100010011111100000001111001111001000",
16#b28# => "1000011100001000100100000000100100111000000011110000001",
16#b23# => "1001010110000000000100000000000001101000011101111001000",
16#b27# => "0001000000111011100100000000001100000000000011111110000",
16#b18# => "0001011100000000000100000000100000011110000001111111000",
16#b2e# => "0000100100001000000100000000000000011010000011110000000",
16#b13# => "1000011110001000100100000000000000000010000011110000000",
16#b22# => "0000111000001000100100000000000001000010000001110000000",
16#b21# => "1001001000001000100100000000000000000010000001110111000",
16#b34# => "0000100010000000100100010011110100000001010001111001000",
16#b19# => "0001101010000000000100000000000010111100000011111110000",
16#b5b# => "1000110010000000100100111100000001000001100011111001000",
16#b56# => "0010110000001100000100000011111100111000011001110100000",
16#b51# => "0010101111111000000100000011111101110100011001110000000",
16#b4d# => "1000110000001000100100111111000001111001111001111001000",
16#b5a# => "0010011000000000100100000011001001101000001011111001010",
16#b54# => "0010101010001000100100000011010000101000001011110000000",
16#b50# => "1010100100001000100100000011100000101000001011110000000",
16#b1b# => "1000110001111000100100010011001100000000101001111001000",
16#b57# => "0010101010001111000100111000000001110101100001111001000",
16#b53# => "1010100101110000100100110100000000110001100001111001000",
16#b4e# => "1010100100000111000100000000000001110000000011111111000",
16#b45# => "0010011011110000000100000000011000101100000011111111000",
16#b4a# => "1010001110000110100100000000011010100100000011111110000",
16#b3d# => "1010010011101000000100000000011001100000000011111110000",
16#b43# => "1001111010000110000100000000000010011100000011111111000",
16#b3b# => "0010000011100000100100000011111100010100011001110000000",
16#b36# => "0001110000001101100100000011111100000100011001111101000",
16#b35# => "0001101100001101000100010011111000011001101000110000000",
16#b2f# => "0001101011010000100100000011111100001100010001110010000",
16#b4c# => "0010011010001000100100000011000100101000010011110000000",
16#b44# => "1010001100001000100100000011001000101000010011110000000",
16#b48# => "1010010100000000100100000001111000000000011001111001000",
16#b3c# => "1010001100001000000100001010110000000001111001111001101",
16#b41# => "0011001000000000100100011100000000101001100001111001000",
16#b3a# => "1001111100001000000100010100000000001101100001111001000",
16#b37# => "0000100010000000100100000000000001000010000001110000000",
16#b4f# => "0010011110001110100100110000000001101101100001111001000",
16#b47# => "1010001101101000100100101100000000100101100001111001000",
16#b49# => "1010010010001000100100000011010001101000010011111000000",
16#b46# => "1001111010001000100100000011100001101000010011111000000",
16#b65# => "0011001100000110100100101000111100010101111001111001000",
16#b3e# => "0001101010001000000100010011111100101000011001111010100",
16#b4b# => "1010010100001110000100100100000001100001100001111001000",
16#b3f# => "1001111001100000100100100000000001011101100001111001000",
16#b64# => "0010000110001000100100000011111100101000011001111100000",
16#b72# => "0001110100000000100100000000000000101010100010000000000",
16#b03# => "0011100000001000000100000000100000010000000000001111000",
16#b6e# => "1000000010001000100100000011011100011111011000000110000",
16#b83# => "1011011110001000000100010110000000101001111001000110000",
16#b82# => "0100000000001011100100100010011000100001111001101100000",
16#b52# => "0100000010001001100100000011111100011000011001111010000",
16#b0a# => "1010100000001000000100010000000000100001111011111001000",
16#b2d# => "0000010100001000000100010110000001011001111011111001100",
16#b85# => "1010111010010101100100000000111001111101100011111001101",
16#bb4# => "1100001101110111100100000001101001011101010001110000100",
16#b5e# => "1101101010001000100100100001101001000001111000001001001",
16#b5d# => "1010111111111111000100101100010001000001100011111001001",
16#b39# => "1010111000111001100100110010110101000001111000001001001",
16#b66# => "0011001100001000100100101111111100101011111000101101000",
16#b42# => "0011001000001000000100101100110101100001100000101001001",
16#b38# => "0010000010001000000100000011111100111100011000101001000",
16#b29# => "0001110110000000000110111000101101000001100011111001001",
16#b84# => "1001010100000000100100110101111001000001111000001001001",
16#bb5# => "1010111010001000000100000000000001000010000001110000000",
16#b87# => "1010111100001000000100000000001100000010000001111110000",
16#bb6# => "1010111010001000000100000000000001000010000001110000000",
16#b5c# => "1011011000001000000100000000111101000010000001110000001",
16#b86# => "1101101111101011100100010100111100100100000000010000101",
16#bb7# => "1100001100001111100100111100001101001101100000011110000",
16#b5f# => "1011011100001000000100000000000001000010000001110000000",
16#af9# => "0111110110001111100100011111111101100011101001111001000",
16#afc# => "0111110110000000100100011111111101110001110001111001000",
16#bb3# => "1111111110000000000110101000101010011101000001110000000",
16#bb2# => "0101100100001000100100011111111101100011110001111001000",
16#b6b# => "0101100110001000000100011111111101111101101001111001000",
16#b6a# => "0011010100001000100100101000001101011100100001111110001",
16#b69# => "1101000100001000000100101011111100100011010001111001000",
16#b68# => "0011010010110000100100101011111101111110101001111001000",
16#b67# => "0011010110000000000100101011111101000001111101111001000",
16#bfc# => "0101100000001000100100000000000001000010000001110000000",
16#ba2# => "0011010110001000000100000001000001011100011001110000000",
16#b7e# => "0100000000000000100100101110010100000001111000101001001",
16#b7b# => "0011111000110000000100000011101000110000011001110000000",
16#b78# => "1011110000001100100100101100101100101101100001011001001",
16#b75# => "1011110110010100100100000010010100110100011001010000000",
16#b76# => "1011101010110000100100101011111100111101111000010000000",
16#afe# => "1011101100001000000110101000101100100001100001000111000",
16#afb# => "1111111100001000000100101010111101011101111001111001001",
16#af8# => "0111110000001000100100000000100011100000000010111111000",
16#afa# => "0111110010000000000100000011010001011111010000000000000",
16#b7c# => "1011110110000000000100000000000001000010000001110000000",
16#b7a# => "1011110010000000000100000010000001110110011001010000000",
16#b79# => "1111111010001000000110000000101011000010000001110000000",
16#b77# => "1011101100001000000100000000000001000010000001110000000",
16#bad# => "1111111010000001000100010011101100100000000110001001000",
16#bae# => "1101011110000011000100110011101000000001111001111001000",
16#bfd# => "1101011110001011000100101111010101110001111001100110000",
16#4ff# => "1111111100000001000100101100010000110000000001110000000",
16#b59# => "0011111000001000100100110110000101110101110011110000001",
16#b74# => "0010110000000000100100000011010000110100001001110000000",
16#b00# => "1011101000000000000100101111010100010101111001111001001",
16#b7d# => "0011111000001000100100000010010100110000011001000000001",
16#b81# => "0011111100011000100100110011101000101101111001100000000",
16#bac# => "1111111100000000100100000000000001000010000001110000000",
16#baf# => "1111111100000000100100000000000001000010000001110000000",
16#4fc# => "1111111000000001000100101100000001000010000001110000000",
16#b7f# => "1011110010001000100100000011111111101110011001010000000",
16#b90# => "1100100100001101000100101111010000100001100110110000000",
16#b8f# => "1100100110011000000100000011001101101100011001110000000",
16#b8c# => "0100011110001010100100011111100100110001111110010000000",
16#b2b# => "0100011100111000000100101111010000011101111110000000000",
16#b88# => "1001010100001010100100011111100001100001111110010000000",
16#b8b# => "1100010100000101100100101110110100011101111110000000001",
16#b55# => "1100010001001000100100101111011001100001111110010101000",
16#baa# => "1111111100000000100110101110010001110001111110001100000",
16#4fd# => "1101011010001000100100100000000101000001100000001001001",
16#b92# => "1100100110011000000100000000000001000010000001110000000",
16#b8e# => "0010101100000000100100000000000001000010000001110110000",
16#b2a# => "1001010010001010100100000000000001000010000001110000000",
16#b94# => "0100110111000000100100011111001000011111101000000000000",
16#b99# => "0100101000001010100100000000100101011000011000000000001",
16#adb# => "1100111110000000000110100111101101011101101001111101000",
16#acb# => "1110110100001000101000000001000000000000000001111111000",
16#b98# => "0110010010001001010010101001000010000000000001110000000",
16#b9c# => "0100110100000101100000000001000001000000000000000000000",
16#b97# => "1100111011000000010000000000000000000000000111110000000",
16#b8d# => "0100101001010000100100000000100100110100000000000000001",
16#b93# => "0100011000000000100100000011001000011100011011110000000",
16#b95# => "0100101000001000100100000011110000011110001000000000000",
16#b96# => "0100101000001000100100000011110000011110001000000000000",
16#b9e# => "0100101010001000100000000000000001000010000001110101000",
16#b9f# => "0101001100001000100000011110101101110101100000001000001",
16#ba5# => "1100111001001000100100000010100100011100011000000000000",
16#ba3# => "0101001100000011110000110011111001100001111000100000001",
16#ba1# => "1101000110001000100100001000110100011101100011110000101",
16#ba0# => "1101000010000000101000000000101100111100011000001010000",
16#b9a# => "1101000000000000010000000011110100011100011000001100001",
16#ba6# => "0100110000001000000000011111110100110100000000000011000",
16#b91# => "0101001110001000000100000001001001011100000001111001001",
16#b9b# => "1100100010000000110000010001100001000001000001111001001",
16#b9d# => "0100110110001000100100000000101101110110000001111000001",
16#ba4# => "0100110010001000100000000000101101110110000001111000001",
16#bb1# => "1100010000001000000000001011111100101001111001110110100",
16#b60# => "1101100010000000101100100101110100100101111001000111001",
16#bb0# => "1011000010000100100000111000010101000001111001110111001",
16#b73# => "0101100010000000000100000001100000011100011000110000001",
16#b71# => "0011100000001000110010000001101101111000000001110000001",
16#b8a# => "0011100110000011101000101001100001000000000110000101001",
16#bf3# => "1100010000001000010000001011001100000000101001110000101",
16#b6f# => "1111100100001000100000000000110100101100000000000000001",
16#ba7# => "1011011110001000110010000010100001000000001001110000001",
16#abf# => "1101110000001011000000101000101101011001100000001001001",
16#b70# => "0011100010001000110010000000101101100110000000010000001",
16#b62# => "0000001110001000100100000000101100000000000010001001001",
16#abc# => "1011000000001000000010011000101100000001100111111100000",
16#abd# => "0101111110000000000100000000000000011100100001110000000",
16#bab# => "0101111010010001000100101000110111011100011000010000001",
16#ba8# => "1011011110000100000000100001101100000001000110101101001",
16#b6c# => "0101010101011101110110001011000101101001101001111010100",
16#b61# => "1011011010000000000100000001101100110000000001001010001",
16#ba9# => "1011011000000100000000100001101100000000100110101011001",
16#b6d# => "1011000010000000100100000000000001000010000001111100000",
16#ab6# => "1101110000001001010100101100000001010100000000000110000",
16#ada# => "1110110100000111000100010110000000101000001000000000100",
16#aca# => "0110010010000111000100010110000000101000001000000000100",
16#ab7# => "1111100110000000000110000000101101000000000000000000000",
16#ad8# => "1110011111011100100000010011111001000001110000001011000",
16#ad9# => "1110110100000000000100100000000000011101100000000000000",
16#ace# => "1110110001110100010110101101000001101101111001000000000",
16#ac8# => "1110011101011100100000000010000001010100000000001010000",
16#ac9# => "0110010010000000000100100000000000011101100000000000000",
16#acc# => "0110010011110100001100111001000001111001111001000000000",
16#ade# => "1110011010000000000100101011001000011000110000111101000",
16#bf0# => "0110111000001101100110000000101010100100000000010000000",
16#bed# => "1110101000001000100110000000101010000000000000001101000",
16#ad7# => "1110011010001000000100010000100111011001110000001110000",
16#acf# => "1110101110110000100100000011001000011100011000000000000",
16#acd# => "1110011000000000000100111100000001111101100001100000000",
16#bf9# => "1111100100000000000100101011000100101001101000110000000",
16#bef# => "1111100010000000000100000000100111111000000000001110000",
16#ad5# => "0111011001011000100110000000101101011000000000000000000",
16#adf# => "1110011000001000000100000011001001010100010000001011000",
16#bf2# => "1111100010000000000100101011001000101001101000110000000",
16#bfa# => "1111100100000000000100101011100000101001101000110000000",
16#bf8# => "0111110110001000000100101011010000101001101000110000000",
16#308# => "1101101000001101100110000000101011000000000000000000000",
16#320# => "0000010000101001100100000000101101111100000000000000001",
16#312# => "1101101010001000000110000000101011111000000111110000000",
16#309# => "0000100010001111100100000011011001011100001000000000000",
16#313# => "0111011100000001000100101011000111011100001000000000000",
16#30a# => "0001000110000000101100000011100101011100011001000000000",
16#321# => "1110101010001000001010000000101100100000000111110100000",
16#f2d# => "1001111110000000000100000000000000111000000000000000000",
16#3cd# => "0001011100000000100110000000111111111100000000010100000",
16#f03# => "1110011010000000100110010111001111010101111000111100000",
16#f16# => "1000000000001000100100000000000000000010000000001010000",
16#f14# => "1000101011011000000100000000100001101100000000001011001",
16#f00# => "1000101110000000000100000011100010010100010000001111000",
16#f05# => "1001111010000000000100011111000111011001001000001110010",
16#f08# => "0000001100000000100000011111001101101001101000100000000",
16#f3c# => "0000010111011101110100101100000001101101100000010000000",
16#f0c# => "0000111010001000100100100111111000000001110011110000000",
16#f09# => "1001111110000000000000011100000000100101100000001011000",
16#f10# => "0000100001011101101000110000000000110001100000010000000",
16#f55# => "0000100110000000010000101000000001011101100000001101000",
16#f20# => "1000000100001000000100000000010000100000011000000000001",
16#f01# => "0001000000000000000100000100000001101001100000000000100",
16#f0d# => "1000011000001000000100000000000101000000000000001110010",
16#f0b# => "1001111000000000000000011100000000110101100000001100000",
16#f11# => "0000100010000000010000100000000001011101100000001011000",
16#f02# => "0010101100000000100100000011001100010110011000000000000",
16#f0e# => "1110000100000001000100101111001000101101101010000000000",
16#f0a# => "1000011011111100000000011100000001110001100000001010000",
16#f13# => "0000100000000000010000000100000000011101100000001100100",
16#f0f# => "1000011110001000100100000000000000000010000000000000000",
16#f21# => "1000000110001011101000110000000000110001100000010000000",
16#f12# => "0001000010000000110000000000010000011100011000001010001",
16#f07# => "1111100000000011100110000100101011101001100000001100000",
16#f06# => "0001101110001001100100100100000010011101100000001111000",
16#f1f# => "0000001000001011100100110111001000000001101000101101000",
16#f18# => "1000110010001000000100101011110000000000101001111001000",
16#f31# => "0010101000001111000100000000000111000000000000001111000",
16#f23# => "1001100100000101100100000000000001000000000000000000000",
16#303# => "0001000110001011100110000000111110101100000000000000000",
16#f19# => "1000000100111000100110011100001110101001100000001011000",
16#f30# => "0110111110001001000100101100000100000000000000001111010",
16#f22# => "1001010110001000100100000011110001101010001000001001000",
16#301# => "0001000000001011100110000000111110111000000000000000000",
16#f1a# => "1000000000000000100110011100001111101001100000000000000",
16#f42# => "1000110010000000100100000011111100110000001000001001000",
16#f33# => "0010000010001000000100110000000001111101100000000000000",
16#f1b# => "1001100010001011100100011100000001101001100000001001000",
16#f28# => "1001100010000101100100000100000000110101100000000000100",
16#f24# => "1001010111010111000100101011100000011101101010100100000",
16#f32# => "1001001101111100000100101000000000000011000000000010000",
16#f29# => "1001100000000101100100101100110001101101101000001110010",
16#f2b# => "1001001110000000000100101111010001101101101010010000000",
16#f26# => "1001010000001000100100000000000001000010000000011001000",
16#f2a# => "1001010100001000100100000011010001101010001000001001000",
16#f3a# => "1001001111010000000100010011101101110101001000000100000",
16#f25# => "0001110100001000000100010011100001000001010000100010000",
16#f27# => "1001010110001000100100000000000001000010000000011001000",
16#a80# => "0101111000001000000100000001000000000010011000000000000",
16#abe# => "0001000010001011100110101111001111101101101010101100000",
16#f2c# => "1010010100001000000100000000101001000000000000001110010",
16#f48# => "0001011010000000000100100000101000101001100000001110000",
16#f3b# => "0001110000101000100100110100011000100101100000001110000",
16#f57# => "0001110000001000100100000000000001000000000000000000000",
16#322# => "1110011110111000100100000000000001000000000000000000000",
16#f3f# => "0101111010001111100010011100101011100101100000001010000",
16#f4a# => "1001111001001000110100110000000001000001100000001001000",
16#f39# => "1010010011000000000100010100000001010101100000000101000",
16#3cf# => "1100010011001000100110000000000101101100000001000000000",
16#323# => "0001000100001000000100000000000000101100000000000000000",
16#f3e# => "0101111100001000000110000000101010100110011000001010000",
16#f3d# => "1001111000001011100000000101000000000001111001111001100",
16#f38# => "0001110000000011100100111001000001000001101000100000100",
16#f04# => "0000001000000000000100000000000000000010000000000000000",
16#340# => "1111010000111001001100101000000011010100000000000000000",
16#17e# => "0011111100001000100100100111001000100101101000110000000",
16#1f9# => "0001000000000000000110000000001001000000000000000000000",
16#18b# => "0000111100001001000100111100010010100100011000001000001",
16#382# => "1100010110000000100110000010000100000000000111110000000",
16#17f# => "1111111111100000000110111100001001011101100000001011000",
16#1f8# => "0011111010001011100100000011000100100100001000000000000",
16#163# => "0111110000000110100000000111100101000001101001110000100",
16#162# => "1100010110000000101000101100000001101101100001010001000",
16#189# => "1011000110001101010110000011010001011100010000000000000",
16#343# => "0100000000001000000100000011001000010110010010000000000",
16#341# => "0010000110111000100100000011100000010100010010000111001",
16#311# => "0010000110000000100100101011100000101001110000000000000",
16#f41# => "1111111110001101000110101100001000101101100000011000000",
16#23e# => "0010000011011101000110000100111110110101100000000000100",
16#2fb# => "1001111010001101101000101100000001101101100000011111000",
16#213# => "0111110010001000110110100011110000011110110000010000000",
16#226# => "0000100110001100100100100011101000110001110000001001000",
16#2fe# => "1001001010001000000000011111011001100001110001001101000",
16#212# => "0111110000001000110110110011111101011110110000000000000",
16#23f# => "1001001100001000000100110011011001100011110001001100000",
16#f43# => "1111111000001000000110111000001000011101100000001010000",
16#2fc# => "0010000000001001000100111111001011101100001000000000000",
16#219# => "1100010111001000100110101100000100110001100001000000000",
16#2ff# => "1000110100000011100000101100000000101101100000010100000",
16#218# => "1111111100001011101111111011111000000001110010100000000",
16#1ab# => "1000110110110000000110111001001000000000101000100000000",
16#f40# => "0101010100001000100110111000000101111001100001010111000",
16#2cf# => "1000110100000000100100010011100001101001010000110000000",
16#21b# => "1110011000001000100100111100000001111101100001100000000",
16#21a# => "1000110111100000100100101011100000101001110000110000000",
16#220# => "0001000110000000000100000000000000000010000000000000000",
16#300# => "1101110110001000100110000000101100110100000000000000000",
16#bc0# => "0110111000001000100100000001111100010100000111110000001",
16#bc1# => "1110000010000000000100000011010001011100001000000000000",
16#bba# => "1110000110000000101000000000011100000000000000001110000",
16#bb8# => "1101110100001000001100000011111111001100000000000000000",
16#bc7# => "1101110010000000000100000001100000111101100010001111100",
16#bc6# => "0110001000001000100100000000101100000100000111110001001",
16#bca# => "0110001000001000000100000001100000010000011000110000001",
16#bc8# => "0110010010001000001000100100100001100101100000000000001",
16#bbb# => "0110010100000000010000000011000101011111001000001110010",
16#bdf# => "0110111110001000100100000000000001100000000010000000000",
16#bc5# => "0101111000001000001000011001000000000001100000001101000",
16#bc4# => "0110001110000000101100000000111001000000000000001000011",
16#bda# => "0110001010000000000100101010101101111101111000000101001",
16#bd9# => "1110110110001101100000000000101101101000000010001100010",
16#bbd# => "1110110000000111100101100011101101001100001010000000001",
16#bc2# => "0101111110000011110000000011010001101101101000000000000",
16#bdc# => "1110000010001101100100100110000000011101111011111001000",
16#bce# => "0110111010001111100100010100101100100110100010000000001",
16#bd8# => "1110110100000000000000000000000000000010000000000000000",
16#bbc# => "0101111010000000000000000000000000000010000000000000000",
16#bcf# => "0110111100001111100100010100101101100110100000000000001",
16#bbf# => "1110011110001101000100100111100000010101110000000000000",
16#b02# => "0101111111100110000100101101101100100011111001111001001",
16#bbe# => "0101111000001111100100100000000001010100000000001111000",
16#bc9# => "0101111000001000000100000011001000100100001000000000000",
16#aea# => "0110010100000001000100101111010001010100001010000000000",
16#bc3# => "1111010100001000000110000000101011100000000111111100000",
16#b04# => "0110111110000000000100000000000001000000000000000000000",
16#380# => "0100000000000000000100000000000000000010000000000000000",
16#302# => "1000000100001000000100000000000000000010000000000000000",
16#bd6# => "1110101010001000000100000000000000000010000000000000000",
16#ae8# => "0110111110001111100010000000101100111100000000001011000",
16#ae7# => "1111010010000000010000000011100000010100010000000000000",
16#be4# => "1111001100001000100010000000101011110100000010000000000",
16#b20# => "1111001011011000001100100111011100110101101001111001000",
16#bdb# => "0110111000001111100100000011011100100100001000000000000",
16#bd5# => "1110110110001000100100010100000001010101100000000000000",
16#b01# => "1110101110110011100100100111100001111101101001111001000",
16#af6# => "1111111110000001000100010011101000100100001000000000000",
16#af5# => "0111101110001000000100000011100000010100010000000000000",
16#bd7# => "0111101100000001000100101011101111110100001000000000000",
16#bb9# => "0110111110001111100100000011011010100100001000000000000",
16#be6# => "1101110110000000101000000011100000010100010000000000000",
16#bd4# => "1110101000000000000100000000000000000010000000000000000",
16#bde# => "0110111000001000000100100101000001000001111011111001000",
16#bd3# => "0110111110001111100100000011010110100100001000000000000",
16#bd2# => "0110100000001000100000000011100000010100010000000000000",
16#b40# => "0110100110001000010000100111011011000001101001111001000",
16#af3# => "1111100110001000100100000000000000000010000000000000000",
16#ae4# => "1111001010000000100111101000000001000001100000010111000",
16#ae3# => "1111001100000000000100010111010110010101101000001010000",
16#30b# => "0111000001011101100110100111101011000001101001111001000",
16#af1# => "1111100100000000100100000000000000000010000000000000000",
16#ae1# => "0111000010001000100100000011100000100100001000001100000",
16#af4# => "1000000100000111000110000000101101101000000010010000000",
16#af0# => "0111101010000000000100000011100000010100010000000000000",
16#ae2# => "1111100110110011100100000011110101110000011000000000000",
16#b80# => "1111001010001000100100100111010110110101101001111001000",
16#ae5# => "1111001100000000100100000000000000000010000000000000000",
16#ae0# => "0111000100001000100100000000110101100100000000011100010",
16#af2# => "1111100100001000000100000000000000000010000000000000000",
16#be5# => "0111000110001011100110000011101011100100001000001101000",
16#be7# => "1111001100000000100100000011110100010100010000000000001",
16#bd0# => "1110110010000000100100000000000000100100000111111111000",
16#bcb# => "0110100010000111100100000011010001011100001000001010000",
16#bcc# => "0110010100001000100100000011010001011000010000001011000",
16#be0# => "1110011010000000000100011100000001000001100011111001000",
16#bcd# => "0111000010000110100100111010000001011110011000000000000",
16#be1# => "1110011100000101000100000011100001010100010000001011000",
16#b10# => "0111000011011000100100100111000101101001101001111001000",
16#bdd# => "0110111000000000100100010000100000010101000010010000001",
16#be3# => "0111000110001000000111000000000011100000000010001111000",
16#be2# => "0111000100001000000100000000000000000010000000000000000",
16#be8# => "0111101000001101100100000000000000000010000001010000000",
16#bfb# => "1111010110000000000100111100000001111101100001100000000",
16#bf5# => "0111110100001000101000111000000000111001100001010000000",
16#bf6# => "0111101100000000101100000000010010011100011000001100001",
16#b63# => "0111110000001000100000111000000000111001100001010000000",
16#bf7# => "1011000010001000101100000000000000000000000000001101000",
16#add# => "1000000011000111100110111100000101111101100001100000000",
16#ad6# => "0110111000000101101000111000000000111001100001010000000",
16#ad4# => "1110101110001000001100000100000000011101100000001100100",
16#adc# => "1110101000001000001100000000010001011100011000001101001",
16#ac7# => "0110001000000101000100110111101100000011111001110010000",
16#ac4# => "0110001101011000000100000000100001010100000010001011001",
16#bf4# => "0110001010000000000110111000101010110001100000000100000",
16#bf1# => "0111101110000000000100111100000001110101110000111010000",
16#ac5# => "1111100010000000100110000100101101011101010001110000100",
16#ad0# => "1111111001111101101001111111000111101111111111111111111",
16#ad1# => "0110100011001101101111111111111110010111010111111111111",
16#ac6# => "0110100011000000100100110011000101100101110000100000000",
16#ab3# => "0110001000001100100100110100000001110101100001100001000",
16#ab4# => "0101100110001100000100110000101101110001100001010000001",
16#aff# => "1101101110000100100100001000000001101010101010111111100",
16#310# => "1111111101011000100110110001101010000011011001000000000",
16#ad2# => "1000000110000000001000000000000100000000000111110000001",
16#ad3# => "0110100001001000010000000000000001010100000000000000000",
16#ab1# => "0110001110001000000100110011111001110001110000100000000",
16#ab2# => "0101100111010000100100011100000001011101000000000000000",
16#ab5# => "1101101100000000000100011111010100011101001000000000000",
16#afd# => "0110111100000001000100101101100101100100011010001110000",
16#ac0# => "1111111011111111111111111111111110111111111111111111111",
16#ac3# => "1111111011111111111111111111111110111111111111111111111",
16#ac1# => "1000000100000000000000000000000001000000000000000000000",
16#ac2# => "1000000100000000000000000000000001000000000000000000000",
16#be9# => "0101111110000000100100000000001000000000000000001111010",
16#bea# => "0101111010000000100100000000010010000000000000001111010",
16#beb# => "0101111100000000100100000000100010000000000000001111010",
16#bee# => "0101111100000000100100000000001101000000000000001110010",
16#bec# => "1110110110000000100100000000000011000000000000001110010",
16#5ec# => "1010001100001001000000000111001000100100001000001010000",
16#31d# => "0101010010001000011001000000100101100100000000010100000",
16#583# => "0111011000000000111001111000001011011101100000001000000",
16#5ed# => "0100000011011000101000000000110001000000000000001010001",
16#571# => "0111011110000101011001111100000111011101100000001011000",
16#3aa# => "0011100011000000100010011101010111000000101000100001000",
16#31f# => "0101010100001000011001000000100101100100000000010100000",
16#5ee# => "1010001010001001000000000111001000100100001000001010000",
16#573# => "0111011000001101001000101011011100101001101000101000000",
16#581# => "0011100010001000111001101011010001011110110000110000000",
16#509# => "1100010010001100100000101100000001101101100010000000000",
16#508# => "0000010000000000110100111100000000000001100001000000000",
16#588# => "0000010110000000000100011111011101011001101000101001000",
16#506# => "1100010110000000000000011100000000111001100000000000000",
16#586# => "0000001000001000010100101111001001101101101010100000000",
16#505# => "1100001110001100000000011100000001111101100000000000000",
16#5ef# => "0000001101111000110100101100000001101101100000010000000",
16#587# => "1100010010000000100100110111011101000001101000101001000",
16#574# => "0001110010001000000100110000000001011001000000010000000",
16#50e# => "1011101001001000000100000000100101100100000010001110000",
16#507# => "1000011100001100000000110111011101011001101000101001000",
16#576# => "1000110000000000100110110100100110011000100000000000000",
16#50f# => "1011101010001011100100000011000101000001101000100000000",
16#577# => "0110100010000011111001000000101111000000000000000000000",
16#50c# => "0011100110001000000100110100000000110100110000110000000",
16#50b# => "1000011000000000000000011100000000000000100000001001000",
16#58a# => "0000010000001000110100011100000001000001100000001001000",
16#58b# => "1100010110000001000000101011011110100100001001001101000",
16#572# => "1100010111001000101100110111011101000001101000101001000",
16#58f# => "1000110001010000100110110100100110000000100000000000000",
16#589# => "0100011101001100000000111000100100111001100000011110000",
16#58e# => "1000110110000000100110110100100110000000100000000000000",
16#512# => "0000111010000000000000111011011101111001101000110000000",
16#544# => "0000100010001011101100111011001001111001101000000000000",
16#526# => "1100010001100001000100101011100111100100001000001101000",
16#513# => "1000110100000000100000011100000001000001100000001001000",
16#58c# => "1000110100000000000000011111100000000000101001110000000",
16#524# => "0100011110000000001100111000000000111001100001010000000",
16#521# => "1000011110000000100000011111011100000000101000101001000",
16#519# => "0001000000000000101100111011001110111001101001110000000",
16#561# => "0100110100000000100100000000100101100100000010001110000",
16#58d# => "1011000010000000100100000000000001011000000000000000000",
16#510# => "1001001001001000001000000000000001000000000000000000000",
16#5cb# => "0000100000000000010110111100000000011101100001100000000",
16#5ad# => "0110010000001000101000101111000100101101101001110000000",
16#522# => "1101011010000000110110111011100000011101101001000000000",
16#50d# => "0001000001001000000100101111011101101101101000110000000",
16#543# => "0001000100001000000000011100000001111101100000000000000",
16#541# => "0010000110001000101100011100000000111001100000000000000",
16#520# => "0010000100000000100100111011001001111001101000110000000",
16#517# => "1100010010001001000000101011100011100100001000001101000",
16#515# => "1100010000000001000000101011010011100100001000001101000",
16#518# => "1000101011100011101100011100000000000000100000000000000",
16#51d# => "1100010110000001000100101011010111100100001000001101000",
16#514# => "0000111110000011100000111011011101111001101000110000000",
16#51e# => "1100010111100001000100101011011011100100001000001101000",
16#51b# => "0000111110001011100000111000000001111001100010000000000",
16#51c# => "1000110000001000101100011100000000000001100000001000000",
16#516# => "0000111100000000000000111011011101111001101000110000000",
16#527# => "1001100010001000100000111011001000111001101010000000000",
16#51f# => "1001001101100000101100011100000000100001100000001001000",
16#591# => "1001010000001000100100011111100000011100110000110000000",
16#52e# => "1100100110000011111001011100101111100101100000000000000",
16#528# => "0001011011001110000000011111011100000000101000100000000",
16#523# => "1001010000000000001100011100000001100101100000001001000",
16#525# => "0001000100001000100000111011000100111001101010000000000",
16#52c# => "1100010000000001000100101000000011100100000000011101000",
16#52d# => "0100011110001001000100101011110111100100001000001101000",
16#590# => "1100010110000001000000101011001011100100001000001101000",
16#592# => "0100110101000111000100100011001101101001101010110000000",
16#596# => "0100101110000000101100100111111100100101101000110000000",
16#52a# => "0100011000001001000100101011111011100100001000001101000",
16#52f# => "1001010100001011100100011100000001100101100000000000000",
16#59b# => "1111010001111000100100011100000000100001100000000000000",
16#59a# => "0100110010001000100100101011010000101001101010100000000",
16#593# => "0100110111000111000100100011001001101001101010110000000",
16#597# => "1100100100001011100100011100000000100000101000001100000",
16#595# => "0100101110001000100000011111110000000000101001110000000",
16#594# => "0100101100000000101100100111011100100101101000110000000",
16#52b# => "0100101011110000001000111011011101111001101010100000000",
16#537# => "1011101000000001001000100000101000000000000000001110000",
16#5e9# => "0001101000001101000100110000000010011101100000001111000",
16#5eb# => "1111010110000000100100101011000100101001101010100000000",
16#59e# => "1100111000000000000000101011000100101001110010100000000",
16#502# => "1100111101111000000100110100000001001110100000000000000",
16#557# => "1000000000001000010110000000000011000000000000001111000",
16#535# => "0001101110001000101000000000110000000000000000001110000",
16#575# => "0001101101001101011001110000100000011101100000000000000",
16#501# => "1011101100000000100000011100000001000001100000001001000",
16#5a1# => "1000000000000000111001000000001111000000000000000000000",
16#59c# => "1101000110000000100000000000000001000000000000000110000",
16#534# => "0001101100001000001000000000110000000000000000001110000",
16#532# => "0001101100001101000100110000000000011101100000000000000",
16#530# => "1000000110000000111001000000001111000000000000001100000",
16#536# => "1101000110000000001000101001110010101001111000101111000",
16#503# => "0001101010001101000100110000000000011101100000000000000",
16#531# => "1000000100001000100100101100000001110101100011010000000",
16#aad# => "0010110000001000100100101111000101101101101001111000000",
16#5f3# => "0001101110001101000100110000000010011101100000001111000",
16#553# => "1111100110001000100100101111000101101101101000110000000",
16#a59# => "1010100110001000101010000000010111000000000000000000000",
16#ab0# => "0010110100000000100100011110000001011101101000110000000",
16#a5b# => "0101100000000000010110000000000001000000000000000000000",
16#aaf# => "0010110110010000101000101111000101101101101001111000000",
16#5fd# => "1011110000000000100000000000000001000000000000000000000",
16#54f# => "1010100000000000000100010011100001101101110010100000000",
16#598# => "0001110100001000000100110000000001011001000000010000000",
16#550# => "1111111010000011010110011100000000100001100000000000000",
16#54e# => "1010100110000000000100010011100001101101110010100000000",
16#53a# => "0010011110111100100100110011111000000001110011110000000",
16#599# => "0001110010001000000100110000000001011001000000010000000",
16#558# => "0010101101100011100100010011100001011000110000110000000",
16#5fe# => "1011110000000000100000000000000001000000000000000000000",
16#546# => "1010100100000000000100110011001001000001010000000000000",
16#54c# => "1010001000001000000100110000100110101111000000011110000",
16#556# => "0110111010000000111001000000101111000000000000000110000",
16#5fc# => "0010110010000000000000011111010001000001101000100000000",
16#547# => "1010100110000000000100000000000000000000000000000001000",
16#54d# => "1010001010001011100100110011100110101111001000001110000",
16#554# => "0110111000001110100100101100000011101101100010001111000",
16#555# => "1001100111111110100100000000000011111100000000001111000",
16#5a8# => "0101010000000001100100110100010101110101100000010000001",
16#5a6# => "0101010010000000000100000000000011000000000000001111000",
16#5a4# => "1100111000100000100100110111100001110101101000000000000",
16#59d# => "0101001000101011000100111011011101111001101000110000000",
16#5a0# => "1100111110100000100100000000000001110100000000000001000",
16#5bc# => "0011100000000001000100101011001110100100010000011101000",
16#5a9# => "1101011010111000000100011000000001110001111010010000000",
16#5a7# => "0101010100000000000100000000000011000000000000001111000",
16#5be# => "0011100010000001000100101011010010100100010000011101000",
16#5ac# => "0101111110000011100100100000101001011101100000001110000",
16#5bf# => "0110010100001000000100000011010011011100001000111111000",
16#5d7# => "1110000110000101000100000000000000000000000010001001000",
16#5b2# => "1110101010001101100000000000000000110000000000001101000",
16#5bd# => "0101100110111000001100111000101011111001100010001111000",
16#5ae# => "0101111101111011100100000000000000011100000000000000000",
16#5d6# => "1110000100000000100100000000000000000000000000001000000",
16#5b7# => "1110000110000000100000000000000001110000000000000000000",
16#5b6# => "1101101000001000101100111011010101111001101001001000000",
16#5b5# => "1101101100001000000000011100000000110101100000000000000",
16#5b4# => "1101101010000000101100111000000001111001100000010000000",
16#5b3# => "1101101000000000000000011100000001100101100000000000000",
16#5b1# => "0101100010001000101100111011010000111001101001110000000",
16#5b0# => "0101100100000000100000011100000000100001100000001100000",
16#605# => "1000101010001101110110101011010001011101101000111010000",
16#604# => "0000001001001000100100011100000000110001100000001000000",
16#606# => "0000001110000000000100101011011000101001110010100000000",
16#5c3# => "0000001111100000000110011000011011000001100000001001000",
16#5c1# => "1110000100100000100100110000010101110001100000010100001",
16#60a# => "0011111010001000100100000011100000000001101000100001000",
16#607# => "0000010100001110000100011011001100000001111000101001000",
16#66b# => "0000010001001000000100011011110000000000101001110000000",
16#60b# => "0011010100001000100100011011100001000001110000101001000",
16#6ae# => "1000011000001000101000101111011101101101101000110000000",
16#60c# => "1101011010001000000000101011001001101001111000110000000",
16#608# => "1000011000000011110110101011010001011101101000111010000",
16#60e# => "0101111000001000000000101111011100101101101001110000000",
16#610# => "1000011100001000001100111000000111111001100000011111000",
16#623# => "0000100101001100100000011100101011110001100001001110000",
16#6c9# => "0001000010001000111001111100100001111101100001100110000",
16#60d# => "0110010100000000101000011000000000000001000000001001000",
16#611# => "0100011010001001000100101011101011100100001000001101000",
16#612# => "1110000010000000100100111011100001111001101001001000000",
16#613# => "0100011100001001000100101011101011100100001000001101000",
16#617# => "1110011010001001000000010100000111110000000000001111000",
16#683# => "1101011000001000100100101011001101101000110000110000000",
16#61e# => "1010001010000000100100110000000000110011100000001001000",
16#60f# => "1000110010000000110110111000101011011101100000001110000",
16#645# => "0100000000001000100100101111000101101101101000110000000",
16#61b# => "0000111011011000001000101111011100101101101010100100000",
16#61a# => "1000110000001000110110111100000000011101100001100000000",
16#619# => "1000110000001000001000101100000001101101100010000000000",
16#618# => "1000110110000000110110111000000000011101100000000000000",
16#616# => "1000110000000000001000101111011101101101101000110000000",
16#676# => "1110000100000000100100111100101000001111000000001110000",
16#615# => "1011101000001000001000010100000001111101100000001010100",
16#609# => "1000101010000000100100000000000110011100000000001111000",
16#61c# => "0000010000000000110110010111001000010101101000110000000",
16#64b# => "1000101111000000000100000011100000110000010000011011000",
16#67f# => "1010010000001101000100011011001001000011110000100010000",
16#54a# => "1010010100001000100100000011010000101000010000110000000",
16#569# => "1010010110001110100100000000000110110100000000001111000",
16#614# => "0011010110000101100010011000010111100001100000000100000",
16#64a# => "1010010101010000100100000000000001000000000000000000000",
16#568# => "1010010100001000000100000000000110110100000000001111000",
16#649# => "1000000000000000000100000000000000000010000000000000000",
16#61f# => "0011100000100010000100000000000000000000000000000010000",
16#61d# => "0000111010001000100100100000000001100001100000010000000",
16#62f# => "0000111000000000100000101011001010101001101010101111000",
16#629# => "0001011001111110110000100000000000100001100011001001000",
16#625# => "0001011001111110110000100000000000100001100011001001000",
16#685# => "0001011001111110110000100000000000100001100011001001000",
16#671# => "0001011111111110110000100000000000100001100011001001000",
16#68b# => "0100011011001000100100110000000000110001100011000111000",
16#688# => "1100010010001100000000100100000000100101100011101001000",
16#62e# => "1100010110000000000000000000100111000000000000001111000",
16#690# => "0011100010100010000100111111001001101001101000111000000",
16#68d# => "1100100011100000000100101011000100111101110000110000000",
16#68a# => "0100011101001000100100110000000001110001100001010110000",
16#62c# => "1100010100000000000100011010000110011101100000001111000",
16#68f# => "0011100100100010000100110100000000110101100101101000000",
16#689# => "0100011001001000100100010011100100011001110010100000000",
16#68c# => "1100010100000000100100100100000000100101100011101001000",
16#62d# => "0100011011010000000000000000000111000000000000001111000",
16#68e# => "0011100010000001000100101011101111100100010000001101000",
16#628# => "1100001110100010000100111100000001111101100001100000000",
16#624# => "1001010010100010000100111000000000111001100001100000000",
16#684# => "1001001010100010000100011100010110011101100001010000001",
16#670# => "1100001000100010000100000000000000111100000001000000000",
16#600# => "0011100010000001000100101011100010100100010000000000000",
16#545# => "0011100000000001000100101011101010100100010000000000000",
16#5a3# => "1010001110000000100100101011010000101001101000110000000",
16#582# => "0011100110000001000100101011100111100100010000001101000",
16#578# => "1000000110000000000100000000000000000010000000000000000",
16#5a2# => "1011110100000011100100000000000001000000000000001111000",
16#580# => "1101000100001011100100000011100001000001101000100000000",
16#5a5# => "0100000111000000000100000011010001000001101000100000000",
16#5e8# => "1000000110001000101010000000000101000000000000000000000",
16#5af# => "1111010010000000000100100000000001011111001000110000000",
16#579# => "1101011000001000111001000000101111100000000000010000000",
16#660# => "1011000111011000101000010011110010111000101000101110000",
16#662# => "1011000000000000011001000000000001000000000010000001000",
16#67d# => "1011000010001101100000101111011101101101101010101010000",
16#67c# => "0011111000000000100000010011100000111000101000101101000",
16#67e# => "0011111110000011111001000000100001000000000000000000000",
16#62b# => "0011111111110000000100000011000101000001101000101100000",
16#627# => "0011111111110000000100000011000101000001101000101100000",
16#687# => "0011111111110000000100000011000101000001101000101100000",
16#673# => "0011111001110000000100000011000101000001101000101100000",
16#661# => "1011000000000000011001000000001101011100000000001011000",
16#62a# => "0101001101111110100100101111011100101101101010101000000",
16#626# => "0101001101111110100100101111011100101101101010101000000",
16#686# => "0101001101111110100100101111011100101101101010101000000",
16#672# => "0101001011111110100100101111011100101101101010101000000",
16#53e# => "1010001100000000000000011111100000000000101001110000000",
16#53c# => "1100010110001001000000101011110011100100001000001101000",
16#539# => "1001111111001000001100111000000000111001100000011000000",
16#6a0# => "0001110010000000100010011100010111111101100000001001000",
16#69f# => "1101000110000000010110000000000001000000000000000000000",
16#693# => "1100111110001000100000011100000000111001100000001001000",
16#692# => "1100100100001000110110101100000000101101100010001000000",
16#695# => "0100101110001000000100011100000000110101100000000101000",
16#694# => "0100101000000000100000111011001001111001101000000000000",
16#6ca# => "0100101110000000001100011100000001110001100000000000000",
16#538# => "0110010100001000000010111000011011111001100010000000000",
16#533# => "0001110110000000001100011100000001100101100000001001000",
16#69c# => "1100010010001001000000101011101111100100001000001101000",
16#6b8# => "0100110011111000000000011111011100000001101000100001000",
16#696# => "1101110111000000001100111011010000111001101001000000000",
16#699# => "1110000110000000110110111000000001011101100000000100000",
16#69e# => "0100110101000000101000101100000001101101100000011010000",
16#69d# => "1100111001001000010110111100000000011101100001100101000",
16#698# => "1100111000000101000100101000000000101000111000110000000",
16#69a# => "0100110110000000000100011111000101011101110010100000000",
16#69b# => "1100010101010000000110111000100001011101100000000100000",
16#6ba# => "0100110100000000000000011111011100000001101000100001000",
16#6a9# => "1101011110000000110110110011100000110001101000110000000",
16#6a3# => "0101010110000000100100110011010000110001101000110000000",
16#63f# => "1101000111100000100000011111000100110001110000110000000",
16#6a4# => "1001111100001000110110101100000001101101100000010000000",
16#6a1# => "0101010001101110000100110011010001110001101000110100000",
16#6a5# => "1001111010001000110110101100000001101101100000010000000",
16#6ad# => "1101011100001000100000011111010001000001101000101001000",
16#6a8# => "1101011000000000110110110011100000110001101000110000000",
16#6aa# => "0101010010000000000000011111000100110001110000110000000",
16#6a6# => "1001111010001000110110101100000001101101100000010000000",
16#632# => "0101010000000000000000110011000100110001110000110000000",
16#637# => "0101010100000000000100110011000100110001110000110000000",
16#634# => "0101010100000000000100110011000100110001110000110000000",
16#633# => "0101010110000000000000110011000100110001110000110000000",
16#620# => "0001110000000000000100101100101010101101100010001110000",
16#636# => "0001000010000000000100101011011101101000110000110000000",
16#630# => "0001101011010000000000000000000001000000000000000000000",
16#635# => "1001100110111101011001000000100001000000000000000000000",
16#6ac# => "0001101011001000100100011000000001011001100000000000000",
16#6a2# => "1101011000000000000100011011001100111101111000101001000",
16#6ab# => "1101000000001000000000011111100000110001101010101001000",
16#6a7# => "0101010000001110010110101100000000101101100000010100000",
16#631# => "0100000000000000100000101111011100101101101000110100000",
16#674# => "0010110110001000101000011000000000100001100000000000000",
16#63a# => "1011101110000000010110000000000001011100000000001000000",
16#650# => "1001111010000011100100101111011101101101101010100000000",
16#63b# => "1010100100000000000100000011000101111101101000100000000",
16#647# => "0001110110001011100000011100000000110101100000000000000",
16#6af# => "1010001010001000111001000011100001000001101000100000000",
16#64c# => "1011110100001000000100000000001011011000000000001111000",
16#64f# => "0010011000000011100100110011100000110001101010100000000",
16#64e# => "0010011011001000100000111000000000000011111010100000000",
16#63c# => "0010011110001000010110000011100000111000010000010000000",
16#64d# => "1011110010001000001000000011001010011000001000001111000",
16#640# => "0010011000000000111001000000001110011100000000000000000",
16#639# => "0001110010000000000100000011100001011100011000010000000",
16#642# => "0001110110000011111001011000001111011101100000001000000",
16#63e# => "0010000101001000001000011000110010000001100000001110000",
16#63d# => "1001111000001000011001000000000011000000000000000000000",
16#638# => "1011110100001000001000000000000111011000000000001111000",
16#6b9# => "1101101000000000110110011100000001111001100001001001000",
16#6b1# => "1101110111000000100000101100000111101101100010001111000",
16#681# => "0101100010000000110110011100101010110001100000001110000",
16#6bc# => "0100011100001001000000101011111010100100010010111101000",
16#6b6# => "0101111001001000001100111000000000111001100000011000000",
16#6b5# => "1101101100001000000000011100000001111101100001101001000",
16#5f8# => "0100011000001001000100101011110111100100010010110000000",
16#6be# => "1100100110000000100000010011010000011001110000110000000",
16#6b4# => "0101111010001000001100111000000001111001100000010000000",
16#6b7# => "1101101110000011100100011100000001111101100000000000000",
16#6b2# => "1101101111001000100000111011011100000001101010001000000",
16#6bb# => "0101100010001000010110011111100000111001101001001001000",
16#5fa# => "1010001110000000000100011111100001000000101001111000000",
16#540# => "0111110001001000000100101111011100101101101001110000000",
16#691# => "0010000100101000000110011100010111110100100000001001000",
16#542# => "0010000110101000000100110100010101110101100000010000001",
16#5cd# => "0110100100000000111001000000101111000000000000000000000",
16#5cf# => "1110011110101000100100110000010100110001100000010000001",
16#55e# => "1010010100000000100000011100000000100001100000000000000",
16#5df# => "1010111100001000011001101100001111101101100000011001000",
16#5f7# => "0110100100000000111001000000101111000000000000000000000",
16#5f9# => "0111110010001000100100100000000001000011111010100010000",
16#559# => "0111110110000000100000011111100001000001101000101001000",
16#5de# => "0010110110000000110110000011100000100000010000010000000",
16#55c# => "1011101110000000100000000000000001111100000000001100000",
16#5f1# => "1010111001001000011001101111001111101101101010011001000",
16#5d3# => "1111100101010000000000110000000001000001111010010000000",
16#5f5# => "0110100110001000110110000000000001000000000000000000000",
16#5fb# => "0111101101111011100100101111010001101101101000110000000",
16#5dd# => "1111010010001000000100011111001000011100110000110000000",
16#5f0# => "0110111010000000111001000000101111000000000000000000000",
16#5f2# => "1111100100000011100100000000000001000000000000000000000",
16#5f4# => "0110100000001000110110000000000001000000000000000000000",
16#a58# => "1101011000001011110110011111001001000001110000101001000",
16#a5a# => "0010110110000101000000100000000001000001111010100000000",
16#aa8# => "0010110100001000010110100011000101100000110000010000000",
16#552# => "0101010000000000000110000000101011000000000000000000000",
16#5f6# => "1010100110001000000100101111010100101101101001110000000",
16#a61# => "1101011101001000101000100000011011100000101001110000000",
16#aae# => "1011000000000000100100100000000000011101111000110000000",
16#5aa# => "0011111110001000100100000000000000011100000000001111000",
16#53d# => "0101010100001101100100000011010001101100010000000110000",
16#53f# => "1001111110100000100100110100010100110101100000011000001",
16#59f# => "1001111110001000100100011000000001100001100000001110000",
16#5ab# => "0000001000000000000100010011000101000001110000101001000",
16#500# => "0011100010000001000100101011011110100100011000001101000",
16#570# => "0011111000000100100100000000000000011100000000000000000",
16#504# => "0011100000000000001000000000000000110100000000001111000",
16#5c7# => "0110010100000000110110000000000001011100000001000000000",
16#5e5# => "0110001100001000101000101100000001101101100010000000000",
16#5c5# => "1111001110000000100100011111110001011101110010100110000",
16#5c8# => "0110001100000000110110000000000001100000000000001000000",
16#5ca# => "0110010110101000000100110100010101110101100000010000001",
16#5c9# => "0000001110000000000100011111100001011101110000110000000",
16#5d1# => "1111010010001000000100011111100000011100110000110000000",
16#5ea# => "1000000100001001001000000100000001000000000000001111000",
16#5d0# => "1111010100001000000100011111010000011100110000110000000",
16#5d4# => "0110100110000000011001000000101111000000000000000000000",
16#67b# => "0011100110000001000100101011010111100100010000001101000",
16#67a# => "1011110000101011000100111100000000111101100000010000000",
16#675# => "1110011000000000101000101100000001101101100000011111000",
16#678# => "1011101111011000110110110000101001011101100000001110000",
16#677# => "1011011010000000000000000000000001000000000000001111000",
16#679# => "1011101001011000110110110000101001011101100000001110000",
16#5d9# => "0011001100001000100100101100000001111001100011011111000",
16#549# => "1110110100000110100100000000000000110100000000000000000",
16#54b# => "1010010010101000100100110100010101110101100000011001001",
16#57c# => "0011001100111000100100010111001000010101101010100000000",
16#57f# => "0011111000000011100100000011010000101100010000000100000",
16#57e# => "0011111110001000100100100011010001011101110001111000000",
16#5d8# => "0011111110111000000100101100000001111001100001001111000",
16#57d# => "1100001010000000000100010111001001010101101010100100000",
16#a67# => "1011011000000000110101100000000000011101100000000000000",
16#a66# => "0011001010001000101000101100000001101101100010001100000",
16#a65# => "0011001110001000010101010000000000011101100000001010000",
16#07d# => "0011001110000001001000101011101010101100010010110000000",
16#081# => "0011111010000000111001101100000100011101100000000000000",
16#011# => "0100000010000000101000000000000001000000000000001111000",
16#010# => "0000100000000000111001010111001000010101101000110000000",
16#a6d# => "0011010101011101101000101100000001101101100010000000000",
16#a68# => "1011011100000000110101100100000001011101100000001101000",
16#a69# => "1011011010000000110101110000000001011101100000001011000",
16#a6b# => "1011011000000000110101110100000000011101100000001100000",
16#a2c# => "0011100000000000000100000000000001101000000000000000000",
16#a64# => "0001011100000000001000010111000100010101101010100000000",
16#a6c# => "0011001110000000010101111100000000011101100000000101000",
16#a6f# => "1011011111011000001000101100000001101101100010000110000",
16#a6a# => "1011011110001000110101101000000000011101100000000000000",
16#a6e# => "1011011100001000110101111000000000011101100000001010000",
16#66a# => "1011011110000000000100000000000001000000000000001111000",
16#668# => "0011010000111000000100101011010001101000101000100111000",
16#669# => "0011100110000001000100101011010111100100010000010000000",
16#657# => "0011100100000001000100101011011111100100010000001101000",
16#658# => "0010101001000001100100100000000000100011100000010000000",
16#6d7# => "0011100010000001000100101011011111100100011000000000000",
16#65a# => "0011010110000011100100000000000011011000000000001111000",
16#654# => "0010110100110000000100000011010001000001101000100101000",
16#a70# => "0010101101000001101010000011011010100000011010111000000",
16#6d6# => "0011100100000001000100101011011111100100011000000000000",
16#6d4# => "1011011110000000100100000000011011011100000000001110000",
16#622# => "1110101110110100100100011100100110101111000000011110000",
16#665# => "0001000110001000001000011111101001000001010000000000000",
16#644# => "0011001110010000111001010000100001011000110000110000000",
16#655# => "1010001110000000000100011000100101011101100000001110000",
16#6d5# => "1110101100000000000100011111100101101111001000110000000",
16#648# => "1110101010000000000100101100000001101101100000010000000",
16#667# => "1010010000000000001000011111011100101101110000100000000",
16#601# => "0110001101011101110110101100000001101101100000010101000",
16#65f# => "1000000110000000100000011111011101011001101010101101000",
16#621# => "1010111010001000100000000011010100101100001010110000000",
16#6c5# => "1000000010000000100000011100000000100101100000001011000",
16#65e# => "1010111100001000100000100111011000101001101000110000000",
16#6bf# => "1010111001011111010110101111001001101101101000000000000",
16#6bd# => "0101111110001000100000011100000001101001100000000000000",
16#66d# => "0101111100000000110110101100101011101101100010001111000",
16#6c7# => "1000000100000000100000011100000000100001100000001100000",
16#65d# => "1010111100001000100100101011010000101001101010100000000",
16#6c6# => "1000000010000000100000011100000000110101100000001010000",
16#65c# => "1010111110001000100000000011000100101000011000010000000",
16#697# => "1110000001000011100100111100000001001111000000000000000",
16#6db# => "0100101010001000100000011111000101000001101000100000000",
16#6b3# => "1110110100001000110110011100000000110001100000000001000",
16#6b0# => "0101100100001000100000101111011101101101101000110000000",
16#6c4# => "0101100100000000000100010100000001111101100000000000100",
16#653# => "1110000011000000100100110100000001110001100000000000000",
16#659# => "1010100110001101001000110100000001110101100010000000000",
16#6c2# => "0010110100000000110110011111000101011101101010100000000",
16#652# => "1010100000001000100100000011111101110100011000010000000",
16#6c0# => "0010110010000000110110011111000101011101101010100000000",
16#6c1# => "0011100000100010001000101111011100101101101000111000000",
16#646# => "1110011100000000100100011111000101011101101000110000000",
16#680# => "1010001000001000010110101111011001101101101010100000000",
16#6cc# => "0100000010000000000000101111011101101101101000110000000",
16#666# => "1110011110001000010110101011010001011101101000110000000",
16#6cd# => "0011001100001000000000000011100001011001101000101001000",
16#6c8# => "1110011100000000100100111000001100011101111000110000001",
16#663# => "0110010010000000010110101100000001101101100000011111000",
16#66e# => "0010000100000000101000000011011000100000001000001110000",
16#664# => "1110110000000000100100000011000100100101110000100010000",
16#66c# => "0011001110000000001000000000011000000000000000001110000",
16#6d2# => "1011011111001000010110110000000000011101100000000000000",
16#6ce# => "0110100101011101101000101100000001101101100000011111000",
16#6d0# => "1110011100001000010110100100000001011101100000001101000",
16#6d1# => "1110011110001000010110100000000001011101100000001011000",
16#6d3# => "1110011000001000010110110100000000011101100000001100000",
16#180# => "1000000010001000100000010111011001010101101010101110000",
16#6e3# => "0100000100000000000110010100000101001100110000000000100",
16#6d9# => "0111000101010111011001000011100100100000011010011010000",
16#6e0# => "0011100100000000000010000000101011011000000000000101000",
16#6dc# => "1000000000001000100000011100000000111101100000001101000",
16#603# => "0110111011011101110101101100000001101101100000010000000",
16#66f# => "1000000110001000100000100011111100101101110000011100000",
16#6e2# => "1011011010001000100100010100011000001100110000001110100",
16#6e1# => "0011100010000000000010100100101011011011100000010101000",
16#6dd# => "1000000110001000100000011100000001111001100000001011000",
16#6df# => "1000000000001000100000011100000001101001100000001100000",
16#6e4# => "1110110010001000000000011100000000110001100000001101000",
16#6da# => "1111001101011101110101101100000001101101100000010000000",
16#6de# => "1110110010001000000000011100000000110101100000001010000",
16#719# => "0011100110000000000110000000101011011000000000000101000",
16#71a# => "1000110110000000100000000000000001000000000000001111000",
16#6e5# => "1110110100001000000000011100000000100101100000001011000",
16#6e7# => "1110110010001000000000011100000000100001100000001100000",
16#71c# => "0000111110000000000011010111001000010101101010100000000",
16#71d# => "0000111100000000011001000000001001000000000000000000000",
16#718# => "0000111100000000100000011100000000101101100000001111000",
16#71b# => "1000110100101000011001000000000101000000000000000000000",
16#6e6# => "1000000000001000000000011100000011011001100000001111000",
16#651# => "1000110000001011100110000000011101000000000000000000000",
16#602# => "1010100000000000100100000011001001000001101000100000000",
16#6f6# => "0111101110000000101000111011011000000001101001110001000",
16#6f5# => "0111101010001101001100111000000001111001100000010000000",
16#6cf# => "0111101110000000101000111000000001111001100000010000000",
16#6cb# => "1110011100001000101100000000000000011100000000000000000",
16#003# => "0110010010001000101010111000011011111001100000010000000",
16#002# => "1000000000001000101100000011001001011100001000110000000",
16#6ec# => "0011100100001000000110000000010110111000000000000000000",
16#6eb# => "0111011110000000001000000000010001110000011000000000001",
16#6ea# => "1111010100001000101100000011011001011100010000000000000",
16#6e9# => "1111010000001000001000000011010000111000001000000001000",
16#6e8# => "1111010110000000101100111011000101011100110000010000000",
16#6d8# => "1111010010000000000100000011010001010100001010000000000",
16#6f7# => "1110110000000000001000000100000001110100100000000000100",
16#682# => "0100000010001000000100000000000001000000000000001111000",
16#641# => "0100000110001000000100010110000001010101111010100000000",
16#643# => "0010000100101000100100000011011001100000001000000000000",
16#6ef# => "0010000000001000100100000000001011000000000000001111000",
16#6ee# => "0111011111001000100100100011110000000001101010101001000",
16#65b# => "0111011000001000000100110100010000000001111001111001001",
16#6fa# => "0111110110101000000100000011001101101100001000000000000",
16#6fe# => "0111110100001000000100000000110100010100000000001101001",
16#6fd# => "1111111000001011100100000000000000110100000000000000000",
16#6ed# => "1111111111001000100100100000000111000001100000001111000",
16#6ff# => "1000000110000000000100000000000000000010000000000000000",
16#6fb# => "1011101000001000101010000000001111110000000000000000000",
16#6fc# => "0111110010001000110100000100011000011100100000001110100",
16#6f9# => "1111111010000000001000101100000001101101100010001111000",
16#6f8# => "0111110000000000110100000000010000011100011000110000001",
16#55d# => "1011110000001000000100100111100001110101110010100000000",
16#5d2# => "1010111111110000100000011111100101100111101010100000000",
16#57b# => "0110100010001000001110000000000000000000000000001101000",
16#51a# => "1011110100001111001000111000000001111001100010000000000",
16#563# => "1000110010001000001110011111100001011101101010100000000",
16#548# => "1011000010001000100000101000000001101001001000110000000",
16#567# => "1010010100000000001110000011010001101100010000001001000",
16#57a# => "1100001100000111000100000000000001011100000000000100000",
16#5dc# => "1011110000001000000100100000000001000001100000001001000",
16#55f# => "0110111010000000000100100111100000110101110000111000000",
16#55a# => "1011000110000000001110000000110001011100000000001110000",
16#562# => "0010110100001110001000000000000001000000000000000000000",
16#551# => "1011000001001000010100100000000000011101100000000000000",
16#5e7# => "1010100110000000101000000011010000101100011000000000000",
16#564# => "1111001100001000110100110111100001011101101010100000000",
16#565# => "0011001010000000001000000011010001101100011000010000000",
16#560# => "1110101010000100101000000011011100110000011000010000000",
16#55b# => "1011000000000000001110000000000000011100000000000000000",
16#5d5# => "1011101000001000100110000000001111110100000000001101000",
16#5e6# => "1100001000000000001000101111011101000000101001110001000",
16#584# => "1111001010001101010100101100000001101101100000010000000",
16#56b# => "1100001100000000110100111011011001111001101000001100000",
16#585# => "0011010100001101101000101100000001101101100000011010000",
16#5e0# => "1111001000000000010100101100000000101101100000011011000",
16#5cc# => "0111000011011101100000000000110000000000000000001110000",
16#56a# => "1110011011001000001110111000000001111001100000010000000",
16#5e4# => "1011011111011101101000000000000001000000000000000000000",
16#5e2# => "1111001110000000010100101111001100101101101000001101000",
16#5ce# => "0111000001011101100000010100000001110011000000000000100",
16#56e# => "1110011100001000001110111011010000111001101010000000000",
16#5e3# => "1111001000000000010100101100000001101101100000011010000",
16#56f# => "1110011110001000001110111000000001111001100000010000000",
16#5e1# => "1111001110000000010100000011010001101100010000001100000",
16#56d# => "1110011100001000001110111011000100111001101010000000000",
16#56c# => "0011001110000000110100110000000000011101100000000000000",
16#a75# => "1011101100001000010100000011100000101100010000010000000",
16#a74# => "1011101010000000100000101111001101101111001000110000000",
16#a73# => "1011101000000000011001000011100010101100001000000010000",
16#a72# => "0011100010001000100100000011001001110100010000110000000",
16#0b0# => "0011100100001000000110001000101010100101100000000100100",
16#a71# => "0011100110001000000100000011010000011000001000000000000",
16#a7a# => "1011110100001000000100110101000001000001111000110000000",
16#a79# => "1011110100001011100100101100000001101101100000011100000",
16#a78# => "1011110110000000101000000011100001000001101000101010000",
16#a77# => "1011110010000000010100100100000000011101100000000000000",
16#a76# => "1011101100001000101000011100101101110001100000000000001",
16#aa5# => "0100000010000000100100110111100001110101101000110000000",
16#a9d# => "1010100100001011111001110000100111011001000000001110000",
16#a8c# => "0100110000001000001000000011010001110100010000110000000",
16#a5c# => "0011111010101000000000011111000101100101010000000000000",
16#a7b# => "1010111010000000010100000000000000100000000001010000000",
16#a7f# => "0011111100001000000000011100000001110001100000000000000",
16#a81# => "0011111010001000111001000000100000011000000011010000000",
16#0ba# => "0101001100000001000100101011001011110100001000110000000",
16#a83# => "1011000000001000100100000000000001011000000000000000000",
16#a98# => "1100111000000011100100000011001000011011101000100000000",
16#a8d# => "0100110111011000001000110011111000000001110011110000000",
16#a7c# => "0100011100000101010100010001101001011100110000111110000",
16#a84# => "0011111110000100100100000000010100100000000000011110000",
16#a86# => "1100001100101011000100100000000001100001100000010000000",
16#a7e# => "1100001110001000000100010000010010011001100000011111000",
16#0b8# => "0101001010000001000100101011000111110100001000110000000",
16#a9c# => "0100000110001011100100110000100101011001000000001110000",
16#a85# => "0011111000000100100100000000010100100000000000011110000",
16#a88# => "1100001110001000000100000000010110000000000000001110000",
16#a63# => "1101110010000000100100110111100001011001101000101001000",
16#a7d# => "0100011010000000100100000000101000000000000000001110000",
16#a8a# => "0011111000000100100100000000010100100000000000011110000",
16#a87# => "1100010011011000000100010000101011011001100000011110000",
16#5c6# => "0101010010000000000100000000000011111100000000001111000",
16#5c4# => "0110001000101000000100100000010100100001100000011101001",
16#5da# => "0110001000000000000100010000110010011001000000001111000",
16#5b9# => "1110110100001101000100110000000001011101100000000111000",
16#566# => "1110011010001000000110000000011011011000000000000000000",
16#50a# => "0011001110001000001000010111001000010101101000110000000",
16#5b8# => "0000010110001000010110100011011001011111001000110000000",
16#53b# => "1101110100000000001000000011001001010000010000110000000",
16#529# => "0001110000001000111001011111100111011101101000000000000",
16#5db# => "1001010010000000100100000011001100011100011000110000000",
16#5ba# => "1101110100101000000100110000010100110001100000010000001",
16#5c2# => "1101110100001000000100000000001011000000000000001111000",
16#5c0# => "1110000110100000000100110000010100110001100000010000001",
16#a8e# => "0100101010001000000100000000000001011000000000000000000",
16#a89# => "0100011000001110000100000011001001110100010000110000000",
16#a92# => "1110011000000000001010000000100000111000000000000000000",
16#a91# => "1110000000000000100110101010011011101000111000110100000",
16#a90# => "1100100010000000101000011111000100100001111000110000000",
16#a99# => "1100100111000000010110000011001001011100001000110000000",
16#a8b# => "0100110010000000100100101111011101101101101010100101000",
16#a8f# => "0100110000001000000100000011001001110100001000110000000",
16#5bb# => "0011001010000000100100010111011000010101101010100000000",
16#a96# => "1101110010001000100010000000010110100000000000000000000",
16#a93# => "1101110010001000100000000000000001001100011000001111000",
16#a9b# => "1100100100001000111001110100100101110111100000000000000",
16#a97# => "1010100100000101100100110000000000011101100000000000000",
16#a94# => "0100101101001000100100000000000001000000000000000000000",
16#aa7# => "0100101000000011100100000011000101000001101000101001000",
16#a54# => "0101001000001000100000011100011000000001100000001110000",
16#a9a# => "0010101010000000011001000000001111100000000000010000000",
16#a51# => "0100000000001000001000010000100100011000110000111110000",
16#aa9# => "1010100110000000111001110000000010011101100000001100000",
16#a55# => "0101010110000000101000000000110010000000000000001110000",
16#a95# => "0010101010000000111001100000001110011111100000001000000",
16#aa4# => "0100000000001000101010000000000011000000000000000000000",
16#a50# => "0101001110000000000100000000000001000000000000001111000",
16#aa2# => "0101010100001000000100010011011101101101010000100000000",
16#a82# => "1101000110111100100100110011100001011111001000110000000",
16#aa6# => "1101110110000101101010101100010111101101100000011100000",
16#aac# => "0101001011010000000100110100000000011101111000111010000",
16#aab# => "1101011000000000010110110111100001110101110000110000000",
16#aaa# => "0101010110001000100100110111010000000001110000100010000",
16#aa3# => "0101010010001000000100010011011101101101010000100000000",
16#a20# => "0100000100001000000100110000000000011001000000000000000",
16#aa1# => "0101010100001000000100011100100111101101100000001110000",
16#a62# => "0001000000000000000100110111001001110101101000110000000",
16#aa0# => "0101010010001000000100011100100110101101000000001110000",
16#a60# => "0100110110001111000100000000000001000000000000000000000",
16#ab9# => "1011000001001000000100000000000001011000000000000000000",
16#88d# => "0100011100001000100100000011001001010000010000000000000",
16#88e# => "0100011000010000100100000000000001000000000000000000000",
16#a30# => "1001111010000110100100011111011101100001110010100000000",
16#88f# => "0110001110000001010110010100000010000000000000001000000",
16#a36# => "0100011010001011100110000100100001011111100000001001000",
16#a32# => "0001101000001011100100011111000101000001110000101001000",
16#a33# => "1001100010000000101000000000000000010000000000000000000",
16#a37# => "0001101001001000000100011111000101000001110000100000000",
16#a2f# => "1001100001111000000100000111000101000001110000100000000",
16#8ea# => "0001011110001000100110000000101010100000000000000000000",
16#8fa# => "1001100101101001011001101000100110011100000000000110000",
16#8ec# => "1000000010000000000000000000000000000010000000000000000",
16#877# => "1111010001010000000000000011100001000001101000100000000",
16#879# => "1011101010001000100100010111001000010101101000110000000",
16#875# => "1011110010000000111001010000100110011011100000000000000",
16#a34# => "1001111000001000000100010111001000010101101010100000000",
16#8ef# => "0111110110001000000100011111011001100001110010100000000",
16#8ed# => "0111011100001110100100100011111101000001110000100000000",
16#8e8# => "0111011100000011100100101000000001101000110000110000000",
16#8ee# => "0100000000000011100100100011001101000001101000100000000",
16#8e9# => "1111001010000101000100000011001001011100001000110000000",
16#a21# => "1111010010000000101010000000100001000000000000000110000",
16#a35# => "0001000010000000110001110100000000011101100000000000000",
16#882# => "0001101100000001000100101011010010110000001000110000000",
16#880# => "0100000110001000000100000011100000110100010000111000000",
16#a48# => "0001101010000101000100000011010001110100010000110000000",
16#a2a# => "0100000000000000000110000000100001000000000000000000000",
16#a47# => "1001010111110000000100100111010001000001110000100000000",
16#a56# => "0100000110000000000110000000100001000000000000000000000",
16#8a1# => "1101000110000000000100100011100001000001101000100000000",
16#a28# => "1111001110001011100110000000100001000000000000000000000",
16#8a0# => "0010101100001011100110010000101010011101100000000000000",
16#881# => "1101000100000011100100100011010001000001101000100000000",
16#a4a# => "0100110100001001000100100011110001010000010000110000000",
16#a46# => "1010010100000100100100000011010000110000001000110000000",
16#a4b# => "1010001111111100000100000100000001011001001000110000000",
16#a25# => "1010010000001000100100100011010000101001101000110000000",
16#a23# => "1010010101000000000100000000000001000000000000000000000",
16#a4c# => "0001000000001011100100000000000001000000000000000000000",
16#a24# => "1010010110001000100100100011010000101001101010100000000",
16#a57# => "1001001100000111000100000000000001000000000000000000000",
16#a22# => "0100110010001001000100100011010101010000010000110000000",
16#a49# => "0010011100000100000100100011100001000001101000100000000",
16#a45# => "1010010100000100100100000011010000110000001000110000000",
16#a4d# => "0100110110001011100110000011100001010000010000110000000",
16#89a# => "0100110100001000100100100111000100100101110000110000000",
16#a44# => "0100101010001001000100100011001101010000010000111010000",
16#891# => "1010111110000000010110111100000000011101100001100000000",
16#87c# => "0011111010001000000100011111000101011101110000110000000",
16#85c# => "1100100000000101101000101100000001101101100010001100000",
16#846# => "1010111010000000010110111011010101011101101001001101000",
16#87e# => "1010001100001000001000000011111100101100011000110000000",
16#883# => "0011111111011000011001000000100111000000000000001010000",
16#897# => "0100000010001000101000111011001101111001101000000000000",
16#89b# => "0100101010001000110001000000000000011100000000001010000",
16#898# => "1010111010001000001100111000000001111001100010001010000",
16#892# => "0100110110000101100100111011011000111001101000001101000",
16#896# => "1100100101011000001000000000000000000000000000001011000",
16#893# => "0100101000001000010110101100000001101101100010000000000",
16#85e# => "1100100110001000100000100011001100100001101010110000000",
16#890# => "1010111100001000001100111000000001111001100010000000000",
16#85d# => "1011101110001001000000011000000011000000000000000000000",
16#894# => "1010111011011000111001000000100110111000000000000000000",
16#8eb# => "0100101000000101101000101100000001101101100010001100000",
16#899# => "1111010000001000110110100001000001011101111000101010000",
16#85f# => "1100001100000000000000011111001001000001110000100000000",
16#895# => "1111010000001000110110000000000000011100000000000101000",
16#a3f# => "1110011010000000100110000000010111000000000000000000000",
16#a40# => "1001111100001110100100010111001000010101101010100000000",
16#a29# => "0010000001101000000100000011010001100000001000110000000",
16#a4f# => "1001010001111000100100000011100001100000010000110000000",
16#a26# => "0010011000001011100100000111010001101001110000110111000",
16#a2e# => "1001001110001100100100011100000001011001100000000000000",
16#a3c# => "0001011110001000000100101011010000101001110000110000000",
16#a2b# => "0001110110001000000100000011001001010000001000110000000",
16#a3e# => "1101000100001000000110000000010111000000000000000000000",
16#a42# => "0001110110001000000100000011001001010000001000110000000",
16#a3b# => "0010000000000000100100000011000101100000010000110000000",
16#a4e# => "0001110011000000100100000011010001101000010000110111000",
16#a27# => "0001110010000101000100011111010101011101110000100111000",
16#a3a# => "0010000110000000100100000011010000101000010000110000000",
16#a43# => "0010000000000000111001000000100110011100000000000000000",
16#a39# => "0010000110001000100100000000000000010000000000000000000",
16#a41# => "1010010010000000101010000000010111000000000000000000000",
16#a38# => "0010000000000000111001000000100111000000000000000000000",
16#a3d# => "0001110000000000100100010111001000010101101010100000000",
16#a31# => "0010000100000000100000101011010001101000110000111001000",
16#8e4# => "1001100000000000100110011100101010100001100000000000000",
16#a9e# => "0100110100001111000100000011010000011000001000110000000",
16#a53# => "1100111010001000000000000011000101010000001000110000000",
16#a9f# => "0100000110001000001000000011001001010000010000110000000",
16#a52# => "1100111000001000100100000011001101011100011000010000000",
16#863# => "0100101100001000100100011111001100011101110000111011000",
16#8e5# => "1011000010001000100100000011001001010000010000110000000",
16#8e7# => "1111001000000101000100000011110001011100001000110110000",
16#8a2# => "0110010010000000100110000000011010000000000000000001000",
16#8b2# => "1101000000001000000100101001000001101000110000110000000",
16#8e6# => "0101100010001000000100111011100001111001101001001000000",
16#8a9# => "1011011000000000000110000000011011000000000000000000000",
16#884# => "0101010000000011100100011100000001111101100000001111000",
16#8b0# => "0001000110000001010110011000011011111000000000001110000",
16#889# => "0101100010000000000100011100100100111101100000001110000",
16#886# => "1100010110000000100100000011011100101100001010110000000",
16#87f# => "1100001110001000000000011111010000101001101000110000000",
16#656# => "0011111011011001011001100000100101011000000000000000000",
16#844# => "0101010000000000000100000011001101010000001000110000000",
16#842# => "0101010100000000000100101111010100111110101000000000000",
16#87d# => "1100001000001000000000011111010000101001101010100000000",
16#845# => "0011100010000001000100101011001011100100010000111101000",
16#843# => "1010001010000011100100000011100100111100010000110000000",
16#878# => "0010000000001011100100000111001001000001101000100000000",
16#876# => "0101010110000000000000011100000001111101100000000000000",
16#8f6# => "1011101000001000011001000000100111000000000000000000000",
16#840# => "1011110110000000001000000111001001000001110000100000000",
16#8bb# => "0010000100000110111001011111100000101111001000010000000",
16#8ae# => "1010010010000000000000000011101001010000001000110000000",
16#8af# => "1101011100001000000100011111010001011101110000110000000",
16#8b1# => "1101011000111000110101101000000001101000110000110000000",
16#8f8# => "0101100010000000100000000011010001101100001000110000000",
16#8f4# => "0111110110000011110110000011111000111100001000110000000",
16#8ac# => "1101011000001000000000111011010001111001101000110000000",
16#8ad# => "1101011011101000000100011111010001011101110000110000000",
16#8f5# => "0111110100000011110110000011011000111100001000110000000",
16#841# => "0111101101101110001000000111010001000001101000100000000",
16#6c3# => "1101110110001001000100100011111000011100010010110000000",
16#8f9# => "0011100100001111000000000000000001111100000000000000000",
16#8f7# => "0111110010000011110110000011011000111100001000110000000",
16#8bc# => "1011011110001000011001000000001111011100000000001011000",
16#8be# => "1101110001111000000100000111001001000001110000101010000",
16#86e# => "0101111111011000001000000000110010000000000000001110000",
16#84d# => "1011011000001000011001000000000011000000000000000000000",
16#84e# => "0010011000000011100100000011111000011100010010111010000",
16#8aa# => "0010011001110000000100000011000101000001101000100000000",
16#872# => "0101010100001110000100011111010000101001101010100000000",
16#84c# => "1101110111111000000100000111001001000001110000100000000",
16#873# => "0101010010001110000100011111010001101001101000111000000",
16#8ba# => "1101101110111011100100000111100001000001110000101100000",
16#8ab# => "1101110010001000000100000111001000000001110000101011000",
16#84b# => "1010010000000000000100000011010101010000001000110000000",
16#8bd# => "1101110100000000100000011100000000000101100000000000000",
16#8c5# => "0101111000111000110000000000000001000000000000000000000",
16#8b8# => "0110001000000100000100000011010000101100001000111000000",
16#84a# => "1010010010000000000100000011000101010000001000110000000",
16#8bf# => "1010010010001110100000111111110000111101101000110000000",
16#8cc# => "1010010000001000100100000011110000111100001000110000000",
16#8b6# => "1110011011011000000100000000000001000000000000000000000",
16#8cb# => "0110001110001110100100000000000001000000000000000000000",
16#8ce# => "1010010010001000100100000011010000111100001000110000000",
16#849# => "0010101010000000100100000000000000000000000000001101000",
16#8ca# => "1110000100001000110101000011000101011100010000110000000",
16#8c9# => "0110010100001011100100000011010000101100001000111101000",
16#8b5# => "0110010010000011100100000111000101000001101000100000000",
16#8f3# => "1010010100000011100100000000000001000000000000001100000",
16#850# => "1111100101011000100000011111001001000001110000100000000",
16#8c8# => "1110011011101000100100000011110100111100001000110000000",
16#8f2# => "1010010110000000000100000011010101010000001000110000000",
16#8f1# => "1110011011101000100100000011010001111100010000111101000",
16#8b4# => "1110011001101000100100000011110000111100001000110000000",
16#8cd# => "1110011010001000100100000011010001111000001000110000000",
16#852# => "1010010010001000100100000011110100111100001000110000000",
16#8cf# => "1111100100001101100100111111100000111101101000110000000",
16#851# => "1110011011101000100000000011110000111100001000110000000",
16#853# => "1010100000000011111001000000100111000000000000000000000",
16#8b7# => "1010100000001011100100000111100001000001101000100000000",
16#8c1# => "1110000010000000000100000011010001111000001000110000000",
16#8c2# => "1110000010000011101000000000000001000000000000000000000",
16#847# => "1110000101001000010000101011001000000001110000101101000",
16#858# => "1010001010001000100000100100000000100101100011101001000",
16#87b# => "0010101100000000100100111100000000011101111000110000000",
16#8a3# => "1011110100001000111001000000100111000000000000000000000",
16#8c0# => "1101000000001000101000000011110000111100001000110000000",
16#85a# => "1010010100000000000000000000000000010000000000000000000",
16#8c3# => "0110001100001110101000000011001000111100001000110000000",
16#85b# => "0010101111001000000100111100000000011101111000110000000",
16#8a6# => "0010110100001000111001100100100110100101100011101001000",
16#8c7# => "0101001110001000000100100000000000100001100011001001000",
16#859# => "0110001100001000100100110100000001110101100001101000000",
16#8b9# => "0010110010000000101000110000000001110001100001010000000",
16#8c6# => "1101110100000000110000011100000000011101100000000000100",
16#89c# => "1100111000001000100100011111010001011101101000110000000",
16#89e# => "1100111110000000010110000000000001000000000000000000000",
16#89d# => "1100111010001101100100000011011100101100001010110000000",
16#89f# => "1011000000001001001000011011011110101100001010111100000",
16#856# => "1100111000001000101000000000000001000000000000001010000",
16#88a# => "0010101010001000010110000000000001111000000000001101000",
16#8e2# => "0111000000000000000100000000000000000000000000000010000",
16#855# => "1100111001101000101000111011100000111001110000111000000",
16#854# => "0010101111100000100000000000000001000000000000001010000",
16#888# => "1100010000001000000100101011000100101001110000110000000",
16#8e0# => "1100100010001000000110000000011011000000000000001100000",
16#8e3# => "0111000010000000000100101011000100000001110000100010000",
16#857# => "0111000110001100000100000011111101101100011000110100000",
16#887# => "0110100100001000000100111011010001111001101000110000000",
16#8f0# => "1100001101100000100100000011011001011100011000010000000",
16#87a# => "1111100110000000000000111000000001111001111000111000000",
16#8fb# => "1011110010001000010110111100000001111101111000110000000",
16#874# => "0111110000001000100000000011011100101100001010110000000",
16#848# => "1011101100000000011001000000100111000000000000000000000",
16#885# => "0110100110001110000100111000000000000001111000101001000",
16#8d2# => "1110110000001000100100111111110001011101101000101000000",
16#8a8# => "0110100110001000000100000011011100101100001010110000000",
16#8d1# => "0100000100000001000100011011111010011100010010110000000",
16#860# => "0110100100000000101000101111011101101101101000110000000",
16#8d0# => "1011000110000011111001000000100110011100000000000000000",
16#862# => "0110100011001000000100111111010001011001101000100000000",
16#8d3# => "1011000010001000000100111111001101000001101000101001000",
16#861# => "1110101010001000100000000000000001000000000000000000000",
16#8e1# => "1110110000000000100000011111010001000001101000100000000",
16#86f# => "0111000100000000110110000000000001000000000000000000000",
16#86d# => "0011010110001000011001000000001110011100000000000000000",
16#8d9# => "1011011110000011100100111111011101011101110010100000000",
16#869# => "1011011000001000101000101100110010101101100000011110000",
16#86b# => "0011010010000000111001110100000010011101100000000000000",
16#8dd# => "0011010100001011100100000011111000110100010010110000000",
16#8dc# => "0110111110000000100100000011000101000001101000100000000",
16#8db# => "0110111000000000000100011111100001000001101001111001000",
16#8d6# => "0011001110000000100100111111010000111101110010100000000",
16#867# => "1110101110001000000100000011001000010000010000111000000",
16#86a# => "0011001001001000101000111111001000111101110000110000000",
16#866# => "1110110100001000001000000000000001010000000000001000000",
16#86c# => "0011001101001000011001000000001111111100000000000000000",
16#865# => "1110101000001000100100111011000100111001110000111011000",
16#8da# => "0011001010000000100100111011100001111001101000110000000",
16#864# => "1110110010001000001000000011010100111100010000110000000",
16#88b# => "0110100000001000100010110100011010110101100000000000000",
16#8b3# => "1100010010001000100100111000000000011101111000111111000",
16#8d8# => "0101100000001000110110101111010000101101101000111000000",
16#868# => "1110110010000000001000000011011100101100001010110000000",
16#8d7# => "0011010100000000011001111100100110011101100000001100000",
16#912# => "1100010110000100000100111011000100011001101000110000100",
16#915# => "0000100101111011000100110000000100011101100000001110010",
16#919# => "1000101000000101100100010011010101011011110000000000000",
16#988# => "1000000010001100100100000000000001110000000000001010000",
16#910# => "1100010100000000000100111011000100011001101000110000100",
16#905# => "0000001111011000000100011100000001110001100000000000000",
16#918# => "0000001010000100000100111000000000011001100000001101100",
16#903# => "1000110111111000000100000000000001000000000000000000000",
16#911# => "0100000110001000000100000011100000000011110001000000000",
16#913# => "0100000000001000000100000011100000000011110001000000000",
16#982# => "0100000110000100111001000000101111000000000000000000000",
16#981# => "0100000010000000100000000000000101000010000000001111010",
16#984# => "1100010010001000000100011111100000011100110000110000000",
16#955# => "1100001110000000011001000000101111000000000000000000000",
16#986# => "1100010100001000000100011111010000011100110000110000000",
16#989# => "1100001101011100111001000000101111000000000000000000000",
16#987# => "1100010010001000000100011111010000011100110000110000000",
16#985# => "1100010100001000000100011111001000011100110000110000000",
16#98a# => "1000000000001000101010000000000101000000000000000000000",
16#980# => "1100010100001000000100011111000100011100110000110000000",
16#904# => "1100001100000000111001000000101111000000000000000000000",
16#9ab# => "1001010000001000000100000011000100011100010000000100000",
16#956# => "1100111110000000100001110000110001011101100000001111110",
16#90d# => "0010101000001000011001000000010110000000000000001011000",
16#957# => "1000011101111100001000000000100101000000000000001110010",
16#900# => "0010101010001101111001000000010111110000000000000000000",
16#929# => "1000000001010000000100110000000000110001100000010110000",
16#9a9# => "1001010110000000100100111011001000000001110000100010100",
16#902# => "0101010100110000100100000000101111000000000000001110010",
16#90e# => "0010101000001000011001000000010111000000000000000000000",
16#90f# => "0000010010001000001000111000110100110001100010001110010",
16#9f0# => "1000011010001000111001111100011011011101100001101011000",
16#917# => "1111100110000000000001000000000001000000000000000111010",
16#916# => "1000101100001000110100000000000001000000000000000000000",
16#92c# => "1000101100001000001000111100000000110101100000000000000",
16#90c# => "0001011110000000011001111011011100011101101001000000000",
16#92f# => "1010111100000000100000000011100001000001101000100000000",
16#9aa# => "1010111110000000100100000011100001000001101000100000000",
16#92d# => "0000111010000000101000110000000000110001100010001001000",
16#91c# => "0001011101001000111001110011011100011101101001011011100",
16#92e# => "0000111011011000000001110011011101000001101000101001100",
16#9a8# => "0001011000001000010000110000000001000001100000001001100",
16#951# => "0000010000001000001000110000000000110101100000000000100",
16#91e# => "1010100010000000111001110000011010011101100001100000100",
16#91d# => "0001011110001000010000110000000001110001100000000000100",
16#953# => "0101010111011000000001110011001001110001101000001000000",
16#930# => "1001100011001000100001110000000000110001100010001010000",
16#9dd# => "1001100110000000010000110011011101000001101000101001100",
16#923# => "0110111100000000100001110011001100110001101000001000010",
16#921# => "0001000010001000110000110000000001000001100000001001100",
16#952# => "0001000100000000100001110011001101110001101000001000000",
16#9dc# => "1010100100001011110000110011111100000001101000100001100",
16#922# => "0110111110000000000001110011100000000000101001110000100",
16#972# => "0001000111001000010000110000110001110001100000011100010",
16#9de# => "1010111110000000100100000011100001000001101000100000000",
16#920# => "0110111001010000000001110011100000000000101001110000100",
16#90a# => "0001000111001000010000110000000000110001100000010000000",
16#938# => "1010111000000000100001000011100001000001101000100000000",
16#939# => "1010111110000000100001000011010001000001101000100000000",
16#933# => "1010111110000000100100000011100001000001101000100000000",
16#935# => "0001110010001000000100000000110000000000000000001100010",
16#93b# => "0001101000000000100001110000110000011101100001001111110",
16#932# => "0001110000110101111001111011010111000011011010000110110",
16#934# => "1001100000001101000001110011111100000001111001101010110",
16#931# => "0001101000111000010000110011111100000001111001001011110",
16#93a# => "0101100110110000000000110011011100110001101010100000000",
16#936# => "0111101010000000100001110011010100110001101001111010010",
16#94d# => "0000010010111101000000011100000001110101100010001001000",
16#945# => "0010011000000000100100011100000001011101100000010000000",
16#944# => "1010001110110000111001111000011010000001100000000001100",
16#941# => "1010001110111000000000011111100000110001101010011001000",
16#940# => "0010000100000000100100011111100001011101101001000010000",
16#93c# => "0010000010000000011001000000011100011000000000000111000",
16#937# => "0011100100001000000001000000110000000000000000001111010",
16#909# => "0001101010001000111001000000010111000000000000000000000",
16#94f# => "0000010100111101000000011100000000110101100000001001000",
16#947# => "0010011010001000100100011100000000011101100001100000000",
16#946# => "1010001000110000111001000000011011000000000000000000000",
16#943# => "1010001100000000000000011111100001110001101010010010000",
16#942# => "0010000110001000100100011111000100011101110001000000000",
16#93e# => "0010000001000000011001000000011100000000000000001000000",
16#908# => "1010010000000000000100111011111101011100111000000000100",
16#948# => "0000010110110000100100011100000001011101100000010000000",
16#90b# => "1010010000110000000100111011111100000000111000000000100",
16#94c# => "1001010000001000000100000011100000011100010000000100000",
16#94e# => "1010010110000000111001110000011011011101100011100000000",
16#949# => "0010011100111000001000000000000001000000000000000110000",
16#94b# => "1010010010000000100100110011111101011101101011000000000",
16#94a# => "1010010101000000111001110011011100011101101011000111000",
16#98c# => "0010110100000000000100000011101101011100010000000011000",
16#997# => "0000111100001000100100111011100000000001110000100010100",
16#98d# => "1101101011011000000100000000110001000000000000001110010",
16#9a7# => "0100011100000011100100000000011001000000000000001110010",
16#99e# => "0101001100001000100100110000000000000001111001111101110",
16#995# => "1100111010110011000100110011010000110001101000000000000",
16#99c# => "0100101110110000100000111011110001000011110000000000100",
16#99d# => "1100111000000000000100010000110011011000100000001100010",
16#9bb# => "1001001110000000100100000011010001101100010000000000000",
16#9ae# => "0000111100001000100100000011011101011100010000000011000",
16#99f# => "0111110110000000000100000000000001000000000000001101010",
16#9b9# => "1111100000001101100100000000000001000000000000000000000",
16#9f7# => "1101110001011000100100000000000000011100000000000000000",
16#9ac# => "0111101010001011100100110011010000110001101000000000000",
16#9f6# => "1101011010110000000100111011010001000001101000100000100",
16#9f8# => "0111101000001000000100000000110011110000000000001110010",
16#9a6# => "0010101010000000100100000000100101000000000000001110010",
16#9a5# => "0101001111010000000100000000000001000000000000000000000",
16#9a3# => "0101001110000101100100000000000101011100000000001111010",
16#9a4# => "1001001000000000100100000011010001101100010000000000000",
16#9a2# => "0101001100000000000100000000000101011100000000001111010",
16#9b7# => "1001010010001000000100000011010100011100010000000100000",
16#9af# => "0000111010001000100100111011100000000001110000100010100",
16#9b3# => "0111110000000000000100000000000001000000000000001101010",
16#97b# => "1111100110001000000100000000000100000000000000001111010",
16#9b5# => "0101111100000011100100110000000000110001100000010000000",
16#9bd# => "1101101110110000100100111011010001000001101000100000100",
16#9b6# => "0101111100000000100100000000101001110000000001001111010",
16#9ad# => "0101100000110011000100010011010000011001101000000000000",
16#9b0# => "1101011100110000100100111011110001000011110000000000100",
16#97a# => "1101000001011011100100111111010000000011000000000010100",
16#9bc# => "1011110000001100100100110000000000011101100000001101110",
16#9b8# => "0101111010000011100001000000000001110000000001001010010",
16#9df# => "1101110000111000010000111011010001000001101000100000100",
16#9f4# => "0110111100001100100001110000000000110001100010001011010",
16#993# => "0111101010000000010000010000101000011000100011011111010",
16#9b1# => "1100100110001011100001110011001101110001101000001001010",
16#9b2# => "0101100110000000110000110000000000000001111001111101110",
16#9ba# => "0101111000001000000001110111000100000001101000101010110",
16#9f5# => "0111101010000000010000110011111100000001111001100110110",
16#992# => "0010110100000000000100000011010001011100010000000011000",
16#9c3# => "0010101010000011100100000000000001000000000000000000000",
16#9bf# => "1110000100001000100100000011100001000001101000101110010",
16#9be# => "1100100110000011100100000000100001000000000000001110010",
16#9c1# => "0101111100001101100100110111000100000001101000101111110",
16#9a1# => "1110000100000011100100000000101001000000000000001110010",
16#9e4# => "1010100010000000000100010000000000011000100000000000000",
16#9c0# => "1111001110000000000100000011011000011100010000000100000",
16#971# => "1001111110001000000100000000000100000000000000001111010",
16#93d# => "0011100000000000100100110000000000011001111000101101110",
16#9c7# => "1001111000000011100100000000110100000000000000001100010",
16#9c6# => "0110001010001000100100110111100001000001101000100000100",
16#990# => "0110001110001000000100000011010000011100010000001100010",
16#9c4# => "1100100100000101000100000000101101000000000000001110010",
16#9c2# => "0110001000000101100100110111000100000001111000100011100",
16#9a0# => "1110000111010000000100000000101001000000000000001110010",
16#954# => "0010101000000000000100000000000001000000000000000000000",
16#9ca# => "0010101110000011100100000000101101000000000000001110010",
16#9c5# => "0110010011010000000100000011100000000011010000100010000",
16#983# => "1111010000001000000100000011010000101100011000000110000",
16#9c8# => "0100000001010000100100000000110011000000000000001110010",
16#978# => "0101111010000000100100000000101000000000000000001111010",
16#9d2# => "0010101010000000100100000000000001000000000000000000000",
16#9d6# => "1001010100001000000100010011111001011101010000110100000",
16#979# => "1000110100001000000100000000000001000000000000000000000",
16#9b4# => "1011110010000101100100000000000001000000000000000000000",
16#9cb# => "1110011100000000100100000000110001000000000000001110010",
16#9d3# => "0110010000001000100100010000010000011000100011011111010",
16#9cc# => "0110100010001101000100000000000001000000000000000000000",
16#9d4# => "1110011111010100100100110000000001110001100010010000000",
16#9ce# => "1110101100110000000100111011001000000001111000100011100",
16#91a# => "1110011000001000000100000000111000110000000001001110010",
16#9c9# => "1110110010000000000100111011000101000011101000100001100",
16#9d1# => "0110010010000000100100000000010011000000000000001110010",
16#9cf# => "0110100110000000100100010011011000011001110000111110010",
16#9cd# => "1110101100110000000100111011000101000011110000100010100",
16#9d0# => "1100100100000000100100000000010011000000000000001110010",
16#9f2# => "0110100100000000000100000000101101000000000000001110010",
16#996# => "1001111110001101101000000000000001000000000000000000000",
16#93f# => "0100101110001000011001110100111010011101100000001100000",
16#994# => "1001111000001000101000110011010001011001110000100000100",
16#98b# => "0100101010111000011001110000111101011101100000001101000",
16#0fd# => "1100010000001001001000100100000110011000000000001111010",
16#00c# => "1111111110000011111001010000110111011101100000001100010",
16#0b7# => "1000011010000000001000110111100001000001101000101101110",
16#00b# => "1101101000001000111001010111010010010101101000110000000",
16#0fc# => "1100010110001001001000100100000110011000000000000111000",
16#998# => "0100110000001000011001011100111101110101100000001101000",
16#99a# => "0100110011011101100000000000000001000000000000000000000",
16#991# => "0100110100001000011001000000111011011000000000000000000",
16#999# => "0100110110001000011001011100110110110001100000001011000",
16#9f1# => "1000000000000000000011010111010000010101101010100000000",
16#99b# => "1111100000000000111001011100010011011001100000000000000",
16#a11# => "1111100010000001011001100100010011000000000000000000000",
16#a03# => "0000100110000000101000000000001000000000000000001111010",
16#a00# => "1000000110001000111001110000010110011101100000000000100",
16#a08# => "1000000000000011100100111011110010000001011010101110110",
16#0c3# => "0000010110000000001010111011101011000001101000101101110",
16#008# => "1110000000001000111001010111010010010101101000110000000",
16#a10# => "1000101100000011000100110000000001011101100000000100100",
16#a0b# => "0000100100000011100100011100000101000001100010001111010",
16#a02# => "0000010100001000100100000011100001000001101000100000000",
16#a01# => "1000000000001011100100111111010000011101100000001110110",
16#009# => "0000010110000000001010111011101011000001101000101101110",
16#a17# => "1111111111001001000100011000100111000000011000001110010",
16#a16# => "1000101100001000100100011111110001110101101010101001000",
16#a14# => "1000101011010000000100111011110101011011110000100010100",
16#a15# => "1000101100000000100100000000000000000010000000000000000",
16#9d9# => "1000000100001000000100000000000000110000000000001011000",
16#9db# => "1110110010000101000100111011001001011001101000100000100",
16#91b# => "1110110010001000100100111011000101000011101000100001100",
16#9d8# => "1001001011001101000100000011010001101100010000000000000",
16#970# => "1110110100000000000000110000000000000001111001111001000",
16#906# => "0011100010000000011001000000010111011000000000011011000",
16#926# => "1100001100000000111001000000101111000000000000000000000",
16#9d5# => "1001001000110000101000101100000001101101100000010000000",
16#925# => "1110101100000000110100101111100101110111010000000000000",
16#9e9# => "1100010000000000101000000011001000011000001000000000000",
16#9ef# => "1111010100000101110100000000100110011000000000011110010",
16#9eb# => "0111011110001000100100111111010000011101100000000000100",
16#9e3# => "1111010100001000101000101100000001101101100000010000000",
16#9ea# => "0111000000111000110100110000000000011101100000000000100",
16#927# => "1111010110001000000100000011010001101100011000000111000",
16#9f3# => "1001001110001000100100000000000001000000000000000000000",
16#9e8# => "1011101110001001001000001111011110110000011000010000000",
16#9e1# => "1111010110001000101000101100000100101101100000011111010",
16#907# => "0011010001010000101000101100000001101101100000010000000",
16#964# => "0000001100001000110100000000000000011100000000000000000",
16#960# => "0011001010000101001000101100000000101101100000010001000",
16#924# => "1011000110000000010100111111001100011101100000000000100",
16#965# => "1011000111011000010100110000000000011101100000000000000",
16#968# => "1011000100000000010100000000000001000000000000000011000",
16#9ec# => "1111010000000000001000000000001100011000000000011110010",
16#9ed# => "0111011111011000010100111100000000011101100001100000000",
16#963# => "0111011110000000101000101100000001101101100010000000000",
16#961# => "1011000000001000110100111000000000011101100001100000000",
16#962# => "1011000100000000101000101111011100101101001000110000000",
16#96b# => "1011000000001000010100111111010001011101100001000000100",
16#9ee# => "1111010110001000001000000011010001101100011010000000000",
16#976# => "0011010100000011100000110111100001000001110001000000100",
16#96a# => "1011101110001000000100110111010001000001110000100000100",
16#9da# => "0011010100001000011001011100011011110001100000000000000",
16#967# => "1110110000001000000000111111001000111001100000000000100",
16#966# => "0011001110001000100100111111000101111101100000000000100",
16#969# => "0011001110001000011001000000011101110100000000001100010",
16#92b# => "0000100010001000100100000000100111000000000000001110010",
16#928# => "1001010110001101100100000011100101011100010000000000000",
16#91f# => "1001010001010000000100000011001100011100010000000100000",
16#901# => "1010111100110000000100000011100000110100010000010000000",
16#950# => "1000000110000000100100000011100001000011110000000000000",
16#973# => "1010100000000000000100000000011001000000000000001110010",
16#92a# => "0011100100001000100100010000111100011000100000001110010",
16#959# => "1001010110001000000100000000010000000000000000001111010",
16#958# => "0010110100000000100100000000110001000000000000001110010",
16#082# => "0011100010001001000100100111010110011000010000001110010",
16#96e# => "1011011000001000100100101111010001101101101010010000000",
16#9d7# => "1011011010001011100100000011100000101100011000011000000",
16#96d# => "1110101100001000100100110111010001000001101000100000100",
16#977# => "1011011010000000100100001000000000011101100000000000100",
16#95c# => "1011101011000000100100000000110011000000000000001110010",
16#96c# => "1011011110000000100100101100000001110001100000000000000",
16#975# => "1011011100000101100100110111010001110101110000000000000",
16#a07# => "1000110000000000100100011100000001011101100000010000000",
16#a0e# => "0000010000000000100100000000101010110100000000001110010",
16#a0a# => "1000011011001101000100110100000000011111100000000111000",
16#974# => "0000010110001000001010101100101011101101100000010000000",
16#96f# => "1011101010000000010100111011010101000001101000101001100",
16#a19# => "1000011100000000000000000000000001000000000000000000000",
16#a05# => "1000110110000011100100110100000001110101100000010000000",
16#a18# => "0000001010110000100100111011010101000001101000100000100",
16#a09# => "1000110110000000000100011111001001011101101000001110010",
16#a0f# => "0000010110000000100100000000101010110100000000001110010",
16#a0d# => "1000011100000000000100011100000001011101100000010000000",
16#a1a# => "1000110000000000111001000000010111000000000000000000000",
16#a1b# => "1000110110001000001000101100000001101101100000010000000",
16#a06# => "1000110010001000100100110100000001011101110000000110000",
16#a0c# => "0000001010111000010100011100000001110101100000001000000",
16#a04# => "0010110100001100101010000000100111110100000000000001000",
16#95b# => "1000011000000001000100000000100111000000000000001110010",
16#9e7# => "1110110110000000000100000000000000011100000000000000000",
16#95a# => "1111001110001101100100101011010100000000101001111001000",
16#9e5# => "1100100000000000100100110000010000101101100000001110010",
16#9e6# => "1111001001011000100100000000000000000000000000001000000",
16#9e2# => "1100100110000000100100000000101101000000000000001110010",
16#95e# => "1010111100001000000100000000000000000010000000000000000",
16#97c# => "1100111000000000000100000000000001000000000000000000000",
16#9e0# => "0011111100000000011001000000010111110000000000000000000",
16#98e# => "0111000110111000000100000011000100011000010000000000000",
16#95f# => "0100011010001101100100000000011011000000000000001110010",
16#95d# => "1010111000001011100100000000000001000000000000001110010",
16#98f# => "1111010000001000000100000011010001101100011000000111000",
-- Replace above this line
others => (others => '0')
);
end package;

package body CCROS is

impure function readCCROS return CCROS_Type is

	variable fileCCROS : CCROS_Type := (others => (others => '0'));
	variable Cline : line;
	variable addr : natural;
	variable CCROSaddr : CCROS_Address_Type;
	file CCROS_lines : text open read_mode is "ccros20130421.txt";

	function fmHex(c : in character) return integer is
	  begin
	  if (c>='0') and (c<='9') then return character'pos(c)-character'pos('0');
	  elsif (c>='A') and (c<='F') then return character'pos(c)-character'pos('A')+10;
	  elsif (c>='a') and (c<='f') then return character'pos(c)-character'pos('a')+10;
	  else 
	  	report "Invalid hex address:" & c severity note;
		return 0;
	  end if;
	  end;

	function fmBin(c : in character) return STD_LOGIC is
	  begin
	  if c='0' then return '0';
	  elsif c='1' then return '1';
	  elsif c='?' then return '0';
	  else
	  	report "Invalid bit:" & c severity note;
		return '0';
	  end if;
	  end;

	-- parity() function returns 1 if the vector has even parity
	function parity(v : STD_LOGIC_VECTOR) return STD_LOGIC is
	variable p : STD_LOGIC;
		begin
			p := '1';
			for i in v'range loop
				p := p xor v(i);
			end loop;
			return p;
		end;
		
	function toString(v : STD_LOGIC_VECTOR) return string is
	variable s : string(1 to 55);
		begin
		for i in v'range loop
			if v(i)='1' then s(i+1):='1';
			else s(i+1):='0'; end if;
		end loop;
		return s;
		end;

	variable char : character;
	variable field : integer;
	variable newC : CCROS_Word_Type;
	variable version : string(1 to 3);
	variable eol : boolean;
	variable cstr3 : string(1 to 3);
	variable cstr8 : string(1 to 8);
	variable cstr55 : string(1 to 55);
	begin
	for i in 1 to 8192 loop
		exit when endfile(CCROS_lines);
		readline(CCROS_lines,Cline);
		exit when endfile(CCROS_lines);
		-- 1-3 = address (hex)
		-- 5-6 = CN hex (ignore 2 lower bits)
		-- 8-11 = CH
		-- 13-16 = CL
		-- 18-20	= CM
		-- 22-23 = CU
		-- 25-28 = CA
		-- 30-31 = CB
		-- 33-36 = CK
		-- 38-41 = CD
		-- 43-45 = CF
		-- 47-48 = CG
		-- 50-51 = CV
		-- 53-55 = CC
		-- 57-60 = CS
		-- 62 = AA
		-- 64 = AS
		-- 66 = AK
		-- 68	= PK
--    File layout:		
--		#AAA  CN CH   CL   CM  CU CA   CB CK   CD   CF  CG CV CC  CS   AAASAKPK

		read(Cline,char);
		if char='#' then next; end if;
		addr := fmHex(char);
		cstr3(1) := char;
		read(Cline,char);	addr := addr*16+fmhex(char);
		cstr3(2) := char;
		read(Cline,char); addr := addr*16+fmhex(char);
		cstr3(3) := char;
		CCROSaddr := CCROS_Address_Type(addr);
--	report "Addr: " & cstr3 severity note;

		-- PN (0) omitted for now
		-- CN
--		read(Cline,char); -- 4
		read(Cline,char); field := fmHex(char);
		read(Cline,char); field := field*16+fmhex(char);
		field := field / 4;
		newC(1 to 6) := conv_std_logic_vector(field,6);
		-- PS (7) and PA (8) omitted for now
		-- CH
--		read(Cline,char);
		read(Cline,char);  newc( 9) := fmBin(char);
		read(Cline,char);  newc(10) := fmBin(char);
		read(Cline,char);  newc(11) := fmBin(char);
		read(Cline,char);  newc(12) := fmBin(char);
		-- CL
--		read(Cline,char);
		read(Cline,char);  newc(13) := fmBin(char);
		read(Cline,char);  newc(14) := fmBin(char);
		read(Cline,char);  newc(15) := fmBin(char);
		read(Cline,char);  newc(16) := fmBin(char);
		-- CM
--		read(Cline,char);
		read(Cline,char);  newc(17) := fmBin(char);
		read(Cline,char);  newc(18) := fmBin(char);
		read(Cline,char);  newc(19) := fmBin(char);
		-- CU
--		read(Cline,char);
		read(Cline,char);  newc(20) := fmBin(char);
		read(Cline,char);  newc(21) := fmBin(char);
 		-- CA
--		read(Cline,char);
		read(Cline,char);  newc(22) := fmBin(char);
		read(Cline,char);  newc(23) := fmBin(char);
		read(Cline,char);  newc(24) := fmBin(char);
		read(Cline,char);  newc(25) := fmBin(char);
 		-- CB
--		read(Cline,char);
		read(Cline,char);  newc(26) := fmBin(char);
		read(Cline,char);  newc(27) := fmBin(char);
  		-- CK
--		read(Cline,char);
		read(Cline,char);  newc(28) := fmBin(char);
		read(Cline,char);  newc(29) := fmBin(char);
		read(Cline,char);  newc(30) := fmBin(char);
		read(Cline,char);  newc(31) := fmBin(char);
		-- PK (32) and PC (33) omitted for now
		-- CD
--		read(Cline,char);
		read(Cline,char);  newc(34) := fmBin(char);
		read(Cline,char);  newc(35) := fmBin(char);
		read(Cline,char);  newc(36) := fmBin(char);
		read(Cline,char);  newc(37) := fmBin(char);
		-- CF
--		read(Cline,char);
		read(Cline,char);  newc(38) := fmBin(char);
		read(Cline,char);  newc(39) := fmBin(char);
		read(Cline,char);  newc(40) := fmBin(char);
		-- CG
--		read(Cline,char);
		read(Cline,char);  newc(41) := fmBin(char);
		read(Cline,char);  newc(42) := fmBin(char);
		-- CV
--		read(Cline,char);
		read(Cline,char);  newc(43) := fmBin(char);
		read(Cline,char);  newc(44) := fmBin(char);
		-- CC
--		read(Cline,char);
		read(Cline,char);  newc(45) := fmBin(char);
		read(Cline,char);  newc(46) := fmBin(char);
		read(Cline,char);  newc(47) := fmBin(char);
		-- CS
--		read(Cline,char);
		read(Cline,char);  newc(48) := fmBin(char);
		read(Cline,char);  newc(49) := fmBin(char);
		read(Cline,char);  newc(50) := fmBin(char);
		read(Cline,char);  newc(51) := fmBin(char);
		-- AA
--		read(Cline,char);
		read(Cline,char);  newc(52) := fmBin(char);
		-- AS
--		read(Cline,char);
		read(Cline,char);  newc(53) := fmBin(char);
		-- AK
--		read(Cline,char);
		read(Cline,char);  newc(54) := fmBin(char);
		-- PK
--		read(Cline,char);
		read(Cline,char);  newc(32) := fmBin(char);
		-- Now fill in PN,PA,PS,PC
		newc(0) := parity(newc(1 to 6)); -- PN = CN
		newc(8) := parity(CONV_STD_LOGIC_VECTOR(CCROSAddr,13)); -- PA = ADDR
--		if (newc(13 to 16)="0010") then
--			newc(32) := parity(newc(22 to 25)); -- PK = CA
--		else
--			newc(32) := parity(newc(28 to 31)); -- PK = CK
--		end if;
		newc(7) := parity(newc(8 to 32) & newc(52) & newc(54)); -- PS = PA CH CL CM CU CA CB CK PK AA AK
		newc(33) := parity(newc(34 to 51) & newc(53)); -- PC = CD CF CG CV CC CS AS

--		Bodge to generate incorrect parity for some locations
		if addr=unsigned'(x"BA0") then -- BA0 has parity change "7" = PS PA PC
--			newc(7) := not newc(7); -- Already doing PA so no need to flip PS
			newc(8) := not newc(8); -- PA
			newc(33) := not newc(33); -- PC
			end if;
		if addr=unsigned'(x"B60") then -- B60 has parity change "B" = PN PA PC
			newc(0) := not newc(0); -- PN
			newc(7) := not newc(7); -- Need to flip PS to keep it correct when PA is flipped
			newc(8) := not newc(8); -- PA
			newc(33) := not newc(33); -- PC
			end if;

		-- Skip over page/location
		read(Cline,char);read(Cline,cstr8);
--		report "Loc: " & cstr8 severity note;
--		for i in newC'range loop
--			if newC(i)='1' then
--				report "1" severity note;
--			else
--				report "0" severity note;
--			end if;
--		end loop;
		-- See if there is a version
		read(Cline,char,eol);
		read(Cline,version,eol);
		if char='-' then
--			report "Version: "&version severity note;
		else
			version := "   ";
		end if;
		
		-- Check for acceptable versions
		-- 000/Blank = Basic
		-- 004 = 64k
		-- 005 = 224UCWs
		-- 006 = Storage Protect
		-- 007 = Decimal Option
		-- 010 = 1050 Console
		-- 014 = Selector Channel #1
		-- 025 = 50Hz timer
		-- A20 = 64k + Storage Protect
		-- Omitted:
		-- 015 = Selector Channel 2
		-- 031 = ??
		-- 906 = Storage Protect Diagnostic
		-- 914 = Selector Channel Diagnostic
		-- 994 = ??
		-- 995 = Local Storage Dump
		-- 996 = Storage Diagnostic
		-- 997 = Mpx Diagnostic
		if version="   " or version="000" or version="004" or version="005" or version="006" or
		version="007" or version="010" or version="014" or version="025" or version="A20" then
			if fileCCROS(CCROSaddr) = (newC'range => '0') then
				fileCCROS(CCROSaddr) := newC;
			else
				report "Duplicate CCROS " & integer'image(CCROSAddr) & " Ver " & version severity note;
			end if;
		else
			report "CCROS " & integer'image(CCROSAddr) & " Ver " & version & " skipped" severity note;
		end if;
--		report "CCROS " & integer'image(CCROSAddr) & ": " & toString(newC);
		end loop;
	return fileCCROS;
	end;

end package body;