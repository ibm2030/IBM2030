---------------------------------------------------------------------------
--    Copyright  2010 Lawrence Wilkinson lawrence@ljw.me.uk
--
--    This file is part of LJW2030, a VHDL implementation of the IBM
--    System/360 Model 30.
--
--    LJW2030 is free software: you can redistribute it and/or modify
--    it under the terms of the GNU General Public License as published by
--    the Free Software Foundation, either version 3 of the License, or
--    (at your option) any later version.
--
--    LJW2030 is distributed in the hope that it will be useful,
--    but WITHOUT ANY WARRANTY; without even the implied warranty of
--    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--    GNU General Public License for more details.
--
--    You should have received a copy of the GNU General Public License
--    along with LJW2030 .  If not, see <http://www.gnu.org/licenses/>.
--
---------------------------------------------------------------------------
--
--    File: ibm2030-vga.vhd
--    Creation Date: 
--    Description:
--    Virtual front panel with indicators via VGA
--    Uses the vga_controller_640-60 module provided by Digilent
--    Page references like "5-01A" refer to the IBM Maintenance Diagram Manual (MDM)
--    for the 360/30 R25-5103-1
--    References like "02AE6" refer to coordinate "E6" on page "5-02A"
--    Logic references like "AB3D5" refer to card "D5" in board "B3" in gate "A"
--    Gate A is the main logic gate, B is the second (optional) logic gate,
--    C is the core storage and X is the CCROS unit
--
--    Revision History:
--    Revision 1.0 2010-07-09
--    Initial Release
--    Revision 1.1 2012-04-07
--		Add Multiplexor Tag indicators
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;

library logic,buses;
use logic.Gates_package.all;
use buses.Buses_package.all;
use work.all;

entity vga_panel IS
	port
	(
		-- Inputs        
		Indicators : in std_logic_vector(IndicatorRange);

		-- Outputs
		Red,Green,Blue,HS,VS : out std_logic;

		-- Clocks
		Clock50 : in std_logic -- 50MHz clock
	);
end entity vga_panel;

architecture behavioural of vga_panel is

-- Layout is 640x480 pixels, divided into 32 columns and 24 rows of 20x20 pixel 'characters'
constant totalLines : integer := 24;
constant totalColumns : integer := 32;
subtype lines is integer range 0 to (totalLines-1);
subtype columns is integer range 0 to (totalColumns-1);
constant totalCharacters : integer := (lines'right+1)*(columns'right+1);
subtype screenCharacterOffset is integer range 0 to totalCharacters-1;

-- Basic screen layout as characters, should correspond to indLayout
type screenType is array(lines,columns) of character;
constant	screen : screenType :=
("    CN   ADR    W         X     ",
 " P012345  P ! P18421  P84218421 ",
 "SA CH   CL    CA  CBCM CU   CK  ",
 " P0123 0123 A0123 0101201AP0123 ",
 "CR  CD        CF  CG CV CC  CS  ",
 " P 0123      012  01 01012A0123 ",
 "           COUNT REG            ",
 "      P84218421 P84218421       ",
 "         DATA    KEY  COMM      ",
 "      P84218421 P8421 8421      ",
 "   FLAGS    TAGS      CHECKS    ",
 "   *****    ****      $$$$$$    ",
 "            *****               ",
 "                                ",
 "    TAGS         BUS OUT        ",
 " stuvwxyz{      P84218421       ",
 "        MSAR         a          ",
 " P84218421 P84218421 b          ",
 "   MSDR       ALU     STAT CHKS ",
 " P84218421 P84218421  cde  fg   ",
 "   B REG     A REG    h i  jkl  ",
 " P84218421 P84218421  mno  pqr  ",
 "A****B****C****D****            ",
 "           F****G****H****J**** "
 );

-- Screen layout in terms of signals, 0 for fixed characters
type screenIndicators is array(lines,columns) of IndicatorRange;
constant indLayout : screenIndicators :=
(
  -- CN,ADRP,W,X
  1=>(1=>1,2=>2,3=>3,4=>4,5=>5,6=>6,7=>7, -- CN
      10=>8, -- PA
		12=>9, -- LP
		14=>10,15=>11,16=>12,17=>13,18=>14,19=>15, -- W
		22=>16,23=>17,24=>18,25=>19,26=>20,27=>21,28=>22,29=>23,30=>24, -- X
		others=>0),
  3=>(1=>25,2=>26,3=>27,4=>28,5=>29, -- SA,CH
      7=>30,8=>31,9=>32,10=>33, -- CL
		12=>34,13=>35,14=>36,15=>37,16=>38, -- AA,CA
		18=>39,19=>40,20=>41,21=>42,22=>43,23=>44,24=>45,25=>46,26=>47,27=>48,28=>49,29=>50,30=>51, -- CB,CM,CU,AK,PK,CK
		others=>0),
  5=>(1=>52, -- PC
      3=>53,4=>54,5=>55,6=>56, -- CD
		13=>57,14=>58,15=>59, -- CF
		18=>60,19=>61, -- CG
		21=>62,22=>63,23=>64,24=>65,25=>66,26=>67,27=>68,28=>69,29=>70,30=>71, -- CV,CC,SA,CS
		others=>0),
  -- Skip SX1 6-12
  -- Skip SX2 13-15
--  13=>(0=>222,1=>218,2=>219,3=>220,4=>221,others => 0), -- P1,2,3,4 for now
--  14=>(1=>223,2=>224,3=>225,4=>226,others => 0), -- T1,2,3,4 for now
--  15=>(0=>235,1=>227,2=>228,3=>229,4=>230,5=>231,6=>232,7=>233,8=>234,others=>0),
  -- End of SX
  15=>(1=>128,2=>129,3=>130,4=>131,5=>132,6=>133,7=>134,8=>135,9=>136, -- Mpx Tags
       16=>137,17=>138,18=>139,19=>140,20=>141,21=>142,22=>143,23=>144,24=>145, -- Mpx Bus
		 others=>0),
  16=>(21=>146, -- MAIN STG
       others=>0),
  17=>(1=>147,2=>148,3=>149,4=>150,5=>151,6=>152,7=>153,8=>154,9=>155, -- M
       11=>156,12=>157,13=>158,14=>159,15=>160,16=>161,17=>162,18=>163,19=>164, -- N
		 21=>165, -- LOC STG
		 others=>0),
  19=>(1=>166,2=>167,3=>168,4=>169,5=>170,6=>171,7=>172,8=>173,9=>174, -- MSDR
       11=>175,12=>176,13=>177,14=>178,15=>179,16=>180,17=>181,18=>182,19=>183, -- ALU
		 22=>184,23=>185,24=>186, -- Stat
		 27=>187,28=>188, -- Chks
		 others=>0),
  20=>(22=>189,24=>190, -- Stat
       27=>191,28=>192,29=>193, -- Chks
		 others=>0),
  21=>(1=>203,2=>204,3=>205,4=>206,5=>207,6=>208,7=>209,8=>210,9=>211, -- B
       11=>194,12=>195,13=>196,14=>197,15=>198,16=>199,17=>200,18=>201,19=>202, -- A
		 22=>212,23=>213,24=>214, -- Stat
		 27=>215,28=>216,29=>217, -- Chks
		 others=>0),
  22=>(1=>218,2=>219,3=>220,4=>221,6=>222,7=>223,8=>224,9=>225,11=>226,12=>227,13=>228,14=>229,16=>230,17=>231,18=>232,19=>233,others=>0),
  23=>(12=>234,13=>235,14=>236,15=>237,17=>238,18=>239,19=>240,20=>241,22=>242,23=>243,24=>244,25=>245,27=>246,28=>247,29=>248,30=>249,others=>0),
  others=>(others => 0));

-- To convert ASCII to the internal 6-bit representation...
-- Not all characters are needed, so some special ones are added
subtype characterCode is std_logic_vector(6 downto 0);
type charArray is array(32 to 123) of characterCode;
constant charTranslate : charArray := (
-- 20->62, 21 ! ->61, 22-23->127, 24->59, 25-29->127, 2A->60, 2B-2F->127
"0111110","0111101","1111111","1111111","0111011","1111111","1111111","1111111",
"1111111","1111111","0111100","1111111","1111111","1111111","1111111","1111111",
-- 30 0 to 39 9 -> 0 to 9, 3A : to 3F ? -> 127
"0000000","0000001","0000010","0000011","0000100","0000101","0000110","0000111",
"0001000","0001001","1111111","1111111","1111111","1111111","1111111","1111111",
-- 40 @ -> 127, 41 A to 4F O -> 10 to 24
"1111111","0001010","0001011","0001100","0001101","0001110","0001111","0010000",
"0010001","0010010","0010011","0010100","0010101","0010110","0010111","0011000",
-- 50 P to 5A Z -> 25 to 35
"0011001","0011010","0011011","0011100","0011101","0011110","0011111","0100000",
"0100001","0100010","0100011",
-- 5B to 60 -> 127
"1111111","1111111","1111111","1111111","1111111","1111111",
-- 61 a to 6F o -> 63 to 77
"0111111","1000000","1000001","1000010","1000011","1000100","1000101","1000110",
"1000111","1001000","1001001","1001010","1001011","1001100","1001101",
-- 70 p to 7A z -> 78 to 88, 7B { -> 89
"1001110","1001111","1010000","1010001","1010010","1010011","1010100","1010101",
"1010110","1010111","1011000","1011001"
);

-- Character bitmaps
-- Fairly self-explanatory
constant characterHeight : integer := 20;
constant characterWidth : integer := 20;
subtype pixLinesRange is integer range 0 to (characterHeight-1);
subtype pixColsRange is integer range 0 to (characterWidth-1);
subtype pixelType is std_logic_vector(1 to 3); -- RGB
subtype pixelRow is std_logic_vector(pixColsRange); -- One scan line
subtype characterRange is integer range 0 to (2**(characterCode'left+1)-1);
type characterGeneratorType is array(characterRange,pixLinesRange) of pixelRow;
constant characterGenerator : characterGeneratorType :=
(	  0 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000111100000000",
			  "00000001111110000000",
			  "00000011100111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011100111000000",
			  "00000001111110000000",
			  "00000000111100000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
     1 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000011000000000",
			  "00000000111000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000111100000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
     2 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000111110000000",
			  "00000001111111000000",
			  "00000011000011000000",
			  "00000000000011000000",
			  "00000000000011000000",
			  "00000000000110000000",
			  "00000000001100000000",
			  "00000000011000000000",
			  "00000000110000000000",
			  "00000001111111000000",
			  "00000011111111000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
     3 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000001111110000000",
			  "00000011111111000000",
			  "00000010000011000000",
			  "00000000000011000000",
			  "00000000000111000000",
			  "00000000011110000000",
			  "00000000000110000000",
			  "00000000000011000000",
			  "00000010000011000000",
			  "00000011111111000000",
			  "00000001111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
     4 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000001100000000",
			  "00000000011100000000",
			  "00000000011100000000",
			  "00000000111100000000",
			  "00000000101100000000",
			  "00000001101100000000",
			  "00000011001100000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000000001100000000",
			  "00000000001100000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
     5 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011111110000000",
			  "00000011111111000000",
			  "00000000000011000000",
			  "00000000000011000000",
			  "00000000000011000000",
			  "00000011111111000000",
			  "00000011111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
     6 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000001111110000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000000000000",
			  "00000011111110000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000001111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
     7 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000000000011000000",
			  "00000000000110000000",
			  "00000000000110000000",
			  "00000000001100000000",
			  "00000000001100000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
     8 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000111100000000",
			  "00000001111110000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000001111110000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000001111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    10 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000011000000000",
			  "00000000111100000000",
			  "00000001100110000000",
			  "00000001100110000000",
			  "00000001000010000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    11 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011111110000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011111110000000",
			  "00000011111110000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000011111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    12 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000001111110000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000001111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    13 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011111110000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000011111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    14 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011111100000000",
			  "00000011111100000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    15 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011111100000000",
			  "00000011111100000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    16 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000001111110000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011001111000000",
			  "00000011001111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000001111111000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    17 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    19 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000000001100000000",
			  "00000000001100000000",
			  "00000000001100000000",
			  "00000000001100000000",
			  "00000000001100000000",
			  "00000011001100000000",
			  "00000011001100000000",
			  "00000011111100000000",
			  "00000001111000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    20=> ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011000011000000",
			  "00000011000110000000",
			  "00000011001100000000",
			  "00000011011000000000",
			  "00000011110000000000",
			  "00000011100000000000",
			  "00000011110000000000",
			  "00000011011000000000",
			  "00000011001100000000",
			  "00000011000110000000",
			  "00000011000011000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    21 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    22 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011000011000000",
			  "00000011100111000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000011011011000000",
			  "00000011011011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    23 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011000011000000",
			  "00000011100011000000",
			  "00000011110011000000",
			  "00000011110011000000",
			  "00000011011011000000",
			  "00000011011011000000",
			  "00000011011011000000",
			  "00000011001111000000",
			  "00000011001111000000",
			  "00000011000111000000",
			  "00000011000011000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    24 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000001111110000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000001111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    25 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011111110000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000011111110000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000011000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    27 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011111110000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000011111110000000",
			  "00000011111000000000",
			  "00000011011100000000",
			  "00000011001110000000",
			  "00000011000111000000",
			  "00000011000011000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    28 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000001111110000000",
			  "00000011111111000000",
			  "00000011000011000000",
			  "00000011100000000000",
			  "00000001110000000000",
			  "00000000111100000000",
			  "00000000001110000000",
			  "00000000000111000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000001111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    29 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011111111000000",
			  "00000011111111000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    30=> ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011111111000000",
			  "00000001111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    31 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011100111000000",
			  "00000011100111000000",
			  "00000001100110000000",
			  "00000001111110000000",
			  "00000000111100000000",
			  "00000000111100000000",
			  "00000000011000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    32 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011011011000000",
			  "00000011011011000000",
			  "00000011111111000000",
			  "00000011100111000000",
			  "00000011000011000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    33 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011100111000000",
			  "00000000111100000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000111100000000",
			  "00000001100110000000",
			  "00000011100111000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    34 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000011000011000000",
			  "00000011000011000000",
			  "00000011100111000000",
			  "00000001111110000000",
			  "00000000111100000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    59 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000001111110000000",
			  "00000011111111000000",
			  "00000111111111100000",
			  "00001111111111110000",
			  "00001111111111110000",
			  "00001111111111110000",
			  "00001111111111110000",
			  "00001111111111110000",
			  "00000111111111100000",
			  "00000011111111000000",
			  "00000001111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    60 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000001111110000000",
			  "00000011111111000000",
			  "00000111111111100000",
			  "00001111111111110000",
			  "00001111111111110000",
			  "00001111111111110000",
			  "00001111111111110000",
			  "00001111111111110000",
			  "00000111111111100000",
			  "00000011111111000000",
			  "00000001111110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    61 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "01100000000111111100",
			  "01100000000111111110",
			  "01100000000110000110",
			  "01100000000110000110",
			  "01100000000111111110",
			  "01100000000111111100",
			  "01100000000110000000",
			  "01100000000110000000",
			  "01100000000110000000",
			  "01111111100110000000",
			  "01111111100110000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    62 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    63 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "10001001000111010001",
			  "11011010100010011001",
			  "10101111110010010101",
			  "10001100010010010011",
			  "10001100010010010001",
			  "00000000000000000000",
			  "01110111110111011110",
			  "10000001001000110001",
			  "01110001001000111110",
			  "00001001001000110010",
			  "01110001000111010001",
			  "00000000000000000000",
			  "00000000000000000000"),
    64 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00001000100010100010",
			  "00010100100010010100",
			  "00111110100010001000",
			  "00100010100010010100",
			  "00100010011100100010",
			  "00000000000000000000",
			  "01110111110111011110",
			  "10000001001000110001",
			  "01110001001000111110",
			  "00001001001000110010",
			  "01110001000111010001",
			  "00000000000000000000",
			  "00000000000000000000"),
    65 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00011111010001000000",
			  "00010000001010000000",
			  "00011100000100000000",
			  "00010000001010000000",
			  "00011111010001000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    66 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "10010110111011010100",
			  "11111001010100110100",
			  "10011111010100011100",
			  "10011001010100110100",
			  "10011001010011010100",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    67 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "01101000100001101001",
			  "10011000100010011001",
			  "11111000100010011001",
			  "10011000100010011111",
			  "10011111111101101001",
			  "00000000000000000000",
			  "10011110010111011110",
			  "10011001010010010000",
			  "10011110010010011100",
			  "11111010010010010000",
			  "10011001010010011110",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    68 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00111111101100111000",
			  "01000001010010100100",
			  "01110001010010111000",
			  "00001001010010101000",
			  "01110001001100100100",
			  "00000000000000000000",
			  "00110111011100000000",
			  "01001100110010000000",
			  "01111100111100000000",
			  "01001100110100000000",
			  "01001111010010000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    69 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00111111101100111000",
			  "01000001010010100100",
			  "01110001010010111000",
			  "00001001010010101000",
			  "01110001001100100100",
			  "00000000000000000000",
			  "01110011001110110000",
			  "01001100100101001000",
			  "01001111100101111000",
			  "01001100100101001000",
			  "01110100101101001000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    70 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00010011001111001100",
			  "00010100101000010010",
			  "00010100101110010010",
			  "00010100100001010010",
			  "00010011001110001100",
			  "00000000000000000000",
			  "00111010010111010010",
			  "00010011010010010010",
			  "00010010110010010010",
			  "00010010010010001100",
			  "00111010010010001100",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    71 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00010011001111001100",
			  "00010100101000010010",
			  "00010100101110010010",
			  "00010100100001010010",
			  "00010011001110001100",
			  "00000000000000000000",
			  "00011100111100110000",
			  "00010010100001001000",
			  "00011100111001001000",
			  "00010100100001011000",
			  "00010010111100111000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    72 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00011100000000000000",
			  "00010010000000000000",
			  "00011100000000000000",
			  "00010010000000000000",
			  "00011100000000000000",
			  "00000000000000000000",
			  "00011100111100110000",
			  "00010010100001000000",
			  "00011100111001011000",
			  "00010100100001001000",
			  "00010010111100110000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    73 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00001100000000000000",
			  "00010010000000000000",
			  "00011110000000000000",
			  "00010010000000000000",
			  "00010010000000000000",
			  "00000000000000000000",
			  "00011100111100110000",
			  "00010010100001000000",
			  "00011100111001011000",
			  "00010100100001001000",
			  "00010010111100110000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    74 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00001100100001001000",
			  "00010010100001001000",
			  "00011110100001001000",
			  "00010010100001001000",
			  "00010010111100110000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    75 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00010010111001001000",
			  "00011110100100111000",
			  "00010010111000110000",
			  "00010010100000110000",
			  "00010010100001001000",
			  "00000000000000000000",
			  "00111010010100101000",
			  "01000010010110101000",
			  "01000011110111101000",
			  "01000010010101101000",
			  "00111010010100101111",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    76 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00001110111101000000",
			  "00010000100001000000",
			  "00001100111001000000",
			  "00000010100001000000",
			  "00011100111101111000",
			  "00000000000000000000",
			  "00111010010100101000",
			  "01000010010110101000",
			  "01000011110111101000",
			  "01000010010101101000",
			  "00111010010100101111",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    77 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00110011010011110000",
			  "01001100111111001000",
			  "01000100110011110000",
			  "01001100110011000000",
			  "00110011010011000000",
			  "00000000000000000000",
			  "01001011011101111000",
			  "01111100110011000000",
			  "01001100110011110000",
			  "01001100110011000000",
			  "01001011011101111000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    78 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "01110001100011100000",
			  "01001010010100000000",
			  "01111010010011000000",
			  "01010010010000100000",
			  "01001001100111000000",
			  "00000000000000000000",
			  "00110111011100000000",
			  "01001100110010000000",
			  "01111100111100000000",
			  "01001100110100000000",
			  "01001111010010000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    79 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "01110001100011100000",
			  "01001010010100000000",
			  "01111010010011000000",
			  "01010010010000100000",
			  "01001001100111000000",
			  "00000000000000000000",
			  "00111001100100000111",
			  "01000010010100001000",
			  "00110011110100000110",
			  "00001010010100000001",
			  "01110011010111101110",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    80 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00111011101110010000",
			  "01000001001001010000",
			  "01000001001110010000",
			  "01000001001010010000",
			  "00111001001001011110",
			  "00000000000000000000",
			  "01110011110011100000",
			  "01001010000100000000",
			  "01110011100101100000",
			  "01010010000100100000",
			  "01001011110011000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    81 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00110011100100101000",
			  "01001010010110101000",
			  "01001011100111101000",
			  "01001010000101101000",
			  "00110010000100101111",
			  "00000000000000000000",
			  "00000011101001000000",
			  "00000001001101000000",
			  "00000001001111000000",
			  "00000001001011000000",
			  "00000011101001000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    82 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00110011100111001110",
			  "01001010010100101001",
			  "01111010010100101110",
			  "01001010010100101010",
			  "01001011100111101001",
			  "00000000000000000000",
			  "00000011101001000000",
			  "00000001001101000000",
			  "00000001001111000000",
			  "00000001001011000000",
			  "00000011101001000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    83 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00111011100110011100",
			  "01000001001001001000",
			  "00110001001111001000",
			  "00001001001001001000",
			  "01110001001001001000",
			  "00000000000000000000",
			  "00000011101001000000",
			  "00000001001101000000",
			  "00000001001111000000",
			  "00000001001011000000",
			  "00000011101001000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    84 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00111011110111001001",
			  "01000010000100101001",
			  "00110011100111001001",
			  "00001010000101000110",
			  "01110011110100100110",
			  "00000000000000000000",
			  "00000011101001000000",
			  "00000001001101000000",
			  "00000001001111000000",
			  "00000001001011000000",
			  "00000011101001000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    85 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00001110111101000000",
			  "00010000100001000000",
			  "00001100111001000000",
			  "00000010100001000000",
			  "00011110111101111000",
			  "00000000000000000000",
			  "00001100100101111100",
			  "00010010100100010000",
			  "00010010100100010000",
			  "00010010100100010000",
			  "00001100111100010000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    86 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00110011100111001110",
			  "01001010010100101001",
			  "01111010010100101110",
			  "01001010010100101010",
			  "01001011100111101001",
			  "00000000000000000000",
			  "00001100100101111100",
			  "00010010100100010000",
			  "00010010100100010000",
			  "00010010100100010000",
			  "00001100111100010000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    87 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00111010010100101110",
			  "01000011110111101001",
			  "01000010010100101001",
			  "01000010010100101001",
			  "00111010010100101110",
			  "00000000000000000000",
			  "00001100100101111100",
			  "00010010100100010000",
			  "00010010100100010000",
			  "00010010100100010000",
			  "00001100111100010000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    88 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00111011110111001001",
			  "01000010000100101001",
			  "00110011100111001001",
			  "00001010000101000110",
			  "01110011110100100110",
			  "00000000000000000000",
			  "00001100100101111100",
			  "00010010100100010000",
			  "00010010100100010000",
			  "00010010100100010000",
			  "00001100111100010000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
    89 => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00111010010111001110",
			  "01000010010100101001",
			  "00110010010111001110",
			  "00001010010100001000",
			  "01110011110100001000",
			  "00000000000000000000",
			  "00001100100101111100",
			  "00010010100100010000",
			  "00010010100100010000",
			  "00010010100100010000",
			  "00001100111100010000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000"),
others => ("00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000111100000000",
			  "00000011111111000000",
			  "00000110000001100000",
			  "00000110000001100000",
			  "00000000000011100000",
			  "00000000000110000000",
			  "00000000001100000000",
			  "00000000011000000000",
			  "00000000011000000000",
			  "00000000000000000000",
			  "00000000011000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000",
			  "00000000000000000000")
);

-- Palette definition
-- Each of the 64 characters has its own palette with a FG and BG
-- colour for the Off and On states
-- The bitmaps above provide the FG/BG selection, the Indicators
-- input signals provide the Off/On selection
subtype sigRange is integer range 0 to 1;
subtype paletteRange is integer range 0 to 1;
type paletteType is array(sigRange,paletteRange) of pixelType;
type fullPaletteType is array(characterRange) of paletteType;
constant characterPalette : fullPaletteType :=
( -- Order is: BGOff FGOff BGOn FGOn
    59 => (("011","000"),("011","100")),-- Chks are red
	 61 => (("011","000"),("011","100")),-- LP is red
	 68 => (("011","000"),("011","100")),-- STOR ADDR is red
	 69 => (("011","000"),("011","100")),-- STOR DATA is red
	 72 => (("011","000"),("011","100")),-- B REG is red
	 73 => (("011","000"),("011","100")),-- A REG is red
	 74 => (("011","000"),("011","100")),-- ALU is red
	 78 => (("011","000"),("011","100")),-- ROS ADR is red
	 79 => (("011","000"),("011","100")),-- ROS SALS is red
	 80 => (("011","000"),("011","100")),-- CTRL REG is red
others => (("011","000"),("011","110"))
);

-- VGA generation
	constant hpixels		: std_logic_vector(9 downto 0) := "1100100000";	 --Value of pixels in a horizontal line (800)
	constant vlines		: std_logic_vector(9 downto 0) := "1000001001";	 --Number of horizontal lines in the display (529)
	
	constant hbp			: std_logic_vector(9 downto 0) := "0010010000";	 --Horizontal back porch (144)
	constant hfp			: std_logic_vector(9 downto 0) := "1100010000";	 --Horizontal front porch (784)
--	constant hbp			: std_logic_vector(9 downto 0) := "0010100000";	 --Horizontal back porch (160)
--	constant hfp			: std_logic_vector(9 downto 0) := "1100000000";	 --Horizontal front porch (768)
	constant	vbp			: std_logic_vector(9 downto 0) := "0000011111";	 --Vertical back porch (31)
	constant vfp			: std_logic_vector(9	downto 0) := "0111111111";	 --Vertical front porch (511)

	signal hc, vc			: std_logic_vector(10 downto 0) := (others=>'0');	 		--These are the Horizontal and Vertical counters
	signal clkdiv			: std_logic := '0';												 	--Clock divider
	signal vidoff			: std_logic;												 			--Tells whether or not its ok to display data
	signal currentLP		: std_logic_vector(5 downto 0) := (others=>'0');			-- Vertical Pixel 0 to 19
	signal currentCP		: std_logic_vector(5 downto 0) := (others=>'0');			-- Horizontal Pixel 0 to 19
	signal currentLine	: std_logic_vector(10 downto 0) := (others=>'0');			-- Line 0 to 23
	signal currentColumn	: std_logic_vector(10 downto 0) := (others=>'0');			-- Column 0 to 31

-- Keyboard handling
	signal keyboard_data_rdy : std_logic;
	signal keyboard_busy : std_logic;
	signal keyboard_error : std_logic;
	
type screenCharacters is array(lines,columns) of characterCode;
-- This function converts the ASCII screen layout into the internal version	
function initScreen (constant screen : screenType) return screenCharacters is
	variable sc : screenCharacters;
	begin
		for r in lines loop
			for c in columns loop
				sc(r,c) := charTranslate(character'pos(screen(r,c)));
			end loop;
		end loop;
		return sc;
	end function;

constant charLayout : screenCharacters := initScreen(screen);


begin
vgaController : entity vga_controller_640_60 port map (
	rst => STD_LOGIC'('0'),
	pixel_clk => clkdiv,
	
	HS => HS,
	VS => VS,
	hcount => hc,
	vcount => vc,
	hchar => currentColumn,
	vchar => currentLine,
	hpixel => currentCP,
	vpixel => currentLP,
	blank => vidoff
	);

	--This cuts the 50Mhz clock in half
	process(Clock50)
		variable currentInd		: IndicatorRange;
		variable currentChar		: characterCode;
		variable pixRow			: pixelRow;
		variable pixPalette		: paletteType;
		variable pix				: pixelType;
		variable fgbg				: paletteRange;
		variable ind				: sigRange;
		begin
			if(Clock50 = '1' and Clock50'EVENT) then
				clkdiv <= not clkdiv;
				currentInd := indLayout(lines(CONV_INTEGER(currentLine)),columns(CONV_INTEGER(currentColumn)));
				currentChar := charLayout(lines(CONV_INTEGER(currentLine)),columns(CONV_INTEGER(currentColumn)));
				if Indicators(currentInd)='1' then ind := 1; else ind := 0; end if;
				pixRow := characterGenerator(characterRange(CONV_INTEGER(currentChar)),pixLinesRange(CONV_INTEGER(currentLP)));
				if pixRow(pixColsRange(CONV_INTEGER(currentCP)))='1' then fgbg := 1; else fgbg := 0; end if;
				pixPalette := characterPalette(characterRange(characterRange(CONV_INTEGER(currentChar))));
				pix := pixPalette(ind,fgbg);
				Red <= pix(1) and not vidoff;
				Green <= pix(2) and not vidoff;
				Blue <= pix(3) and not vidoff;
			end if;
	end process;

END behavioural; 
